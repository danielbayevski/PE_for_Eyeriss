`include "Eyeriss_Row_PE.v"
`include "clock.sv"
`include "FIFObuffer16b_16b.v"
module Eyeriss_Row_tb();


parameter ARRAY_ROW_NUM=2;
reg [18:0] dismod;
reg clrr;
reg [15:0] filterp,mapp;
reg [31:0] pp;
reg [7:0] idp;
reg gm, gf, gp;
wire [15:0] filter,map;
clock clk(.CLK(CLK));
wire [31:0] out, done;
reg start;
reg [3:0]maplen;
reg [7:0] fillen;

wire getdata_fil,getdata_map,getdata_psum;
reg [31:0] expctdoutput [11:0];
wire [15:0] psum_out;
wire pnm;
wire  [51:0] conf;
wire [58:0] GLB_BUS;
wire read;


Eyeriss_Row_PE Row (
 .GLB_BUS(GLB_BUS),
.CLK(CLK),.clr(clrr),
.conf(conf),
.stall(1'b0),
.read(read),
.psum_out(psum_out),
.ready_for_input(), .output_ready(pnm) //empty to front, full to back 
);




//wire getdata_fil,getdata_map,getdata_psum;
//wire [15:0] map, filter;
wire [7:0] id;
wire [31:0] psum_from_PE [2:0];
wire [15:0] Psum_from_GLB;
wire psum_full[2:0] , psum_empty[2:0];
assign GLB_BUS={                          //GBL BUS 		 74 bits
	getdata_fil,           //gather filter to fifo   1  bit
	getdata_map,           //gather map  to fifo     1  bit
	getdata_psum,          //gather GLB PSUM to fifo 1  bit
	map,	        	   //map data to fifo        16 bits
	filter,	        	   //map filter to fifo      16 bits
	id, 	        	   	   //current PE_unit ID      8  bits
	Psum_from_GLB	 	   //PSUM data to fifo       16 bits
    };

/*
Eyeriss_PE pe(.map(map), .filter(filter),.Psum_from_GLB(p),.Psum_from_PE(16'b0),.getdata_fil(gf),.getdata_map(gm),.getdata_psum(gp),
.id_in(8'b1),.stall(1'b0),.psum_i_empty(1'b0),.psum_i_full(1'b0),
 
.CLK(CLK),
.clr(clr),
.conf_i({6'b110000,maplen,fillen,8'b00000001}),
							// enable, GLB input, 0 mult bit, 4 map len,7 fitler len, id =1; 
							//	1bit	1bit 	   4bit			4bit		8bit		8bit 
.ready(),.psum_out(psum_out),.psum_o_empty(pnm),.psum_o_full(),.start(start)
);
*/
/*        conf_i = 
  wire conf_enable;                                               1
	wire conf_psum_input;  //0- psum from PE, 1-psum from GLB     1
    wire [3:0]mult_bit_select;                                    0000
	wire [3:0] conf_maplen;                                       0010
    wire [7:0] conf_filterlen;                                    00000011
	wire [7:0] conf_id;                                           00000001
	=> 11000000100000001100000001
*/     


reg rid,pnd,png;
reg[15:0]check0,chkreg,chkreg2,chkreg3;
wire [15:0] outcheck0;
assign clr=clrr;
assign filter=filterp;
assign map=mapp;
assign Psum_from_GLB=pp;
initial rid=0;
initial check0=0;
assign id=idp;
assign getdata_fil=gf;
assign getdata_map=gm;
assign getdata_psum=gp;



FIFObuffer16b_16b Fifo_outside(
.Clk(CLK),
.dataIn(chkreg),
.RD(rid),
.WR(!pnd),
.EN(1'b1),
.dataOut(outcheck0),
.Rst(clrr),.EMPTY(),
.FULL(read)
);


/*
assign conf[9]={6'b100000,maplen,fillen,8'b00001001};
assign conf[8]={6'b100000,maplen,fillen,8'b00001000};
assign conf[7]={6'b100000,maplen,fillen,8'b00000111};
assign conf[6]={6'b100000,maplen,fillen,8'b00000110};
assign conf[5]={6'b100000,maplen,fillen,8'b00000101};
assign conf[4]={6'b100000,maplen,fillen,8'b00000100};
assign conf[3]={6'b100000,maplen,fillen,8'b00000011};
assign conf[2]={6'b100000,maplen,fillen,8'b00000010};*/
assign conf[51:26]={6'b100000,maplen,fillen,8'b00000001};
assign conf[25:0]={6'b110000,maplen,fillen,8'b00000000};
 initial dismod=0;
always@(posedge CLK) begin
 dismod<=dismod+1;
 pnd<=pnm;
 png<=pnd;
 chkreg<=psum_out;
 chkreg2<=chkreg;
 chkreg3<=chkreg2;
 
 case(dismod)
/* 
 default: 
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
   clrr<=0;
   filterp<=0;
   mapp<=0;
   
   end 
 */
//XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX




19'd0: begin  
  clrr<=1;
 end   
19'd1: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=45;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=21977;
 end   
19'd2: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=81;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=23436;
 end   
19'd3: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=27;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd4: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=61;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd5: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=91;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd6: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=95;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd7: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=42;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd8: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=27;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd9: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=36;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd10: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=91;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd11: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=47;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=41565;
 end   
19'd12: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=26;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=45579;
 end   
19'd13: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=71;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd14: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=38;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd15: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=69;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd16: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=12;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd17: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=67;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd18: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=99;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd19: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=35;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd20: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=94;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd21: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd163: begin  
rid<=1;
end
19'd164: begin  
end
19'd165: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd166: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd167: begin  
rid<=0;
end
19'd301: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=11;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11767;
 end   
19'd302: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=53;
   mapp<=33;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12209;
 end   
19'd303: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=68;
   mapp<=73;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12584;
 end   
19'd304: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=47;
   mapp<=64;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=12207;
 end   
19'd305: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=44;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd306: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd307: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=57;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd308: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd309: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=16;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=25288;
 end   
19'd310: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=35;
   mapp<=23;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=21086;
 end   
19'd311: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=90;
   mapp<=41;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=25762;
 end   
19'd312: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=42;
   mapp<=29;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=21391;
 end   
19'd313: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=88;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd314: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=6;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd315: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=40;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd316: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=42;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd317: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd459: begin  
rid<=1;
end
19'd460: begin  
end
19'd461: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd462: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd463: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd464: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd465: begin  
rid<=0;
end
19'd601: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=70;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4039;
 end   
19'd602: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=50;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5127;
 end   
19'd603: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=6;
   mapp<=90;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10063;
 end   
19'd604: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=1;
   mapp<=29;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5702;
 end   
19'd605: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=93;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=7835;
 end   
19'd606: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=48;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6909;
 end   
19'd607: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=29;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=10635;
 end   
19'd608: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=23;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=8032;
 end   
19'd609: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=84;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd610: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=54;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd611: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=56;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd612: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=8;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=11033;
 end   
19'd613: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=44;
   mapp<=66;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12150;
 end   
19'd614: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=39;
   mapp<=76;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=16234;
 end   
19'd615: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=26;
   mapp<=31;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=12250;
 end   
19'd616: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=23;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=14643;
 end   
19'd617: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=37;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=14807;
 end   
19'd618: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=38;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=20474;
 end   
19'd619: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=18;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=17639;
 end   
19'd620: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=82;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd621: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=29;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd622: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=41;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd623: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd765: begin  
rid<=1;
end
19'd766: begin  
end
19'd767: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd768: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd769: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd770: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd771: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd772: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd773: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd774: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd775: begin  
rid<=0;
end
19'd901: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=6;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8907;
 end   
19'd902: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=73;
   mapp<=58;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11127;
 end   
19'd903: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=86;
   mapp<=4;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11036;
 end   
19'd904: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=21;
   mapp<=30;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=11105;
 end   
19'd905: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=45;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd906: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=24;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd907: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=72;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd908: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd909: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=86;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=26936;
 end   
19'd910: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=90;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=27201;
 end   
19'd911: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=61;
   mapp<=73;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=26751;
 end   
19'd912: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=36;
   mapp<=97;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=27498;
 end   
19'd913: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=55;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd914: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=67;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd915: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=55;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd916: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=74;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd917: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd1059: begin  
rid<=1;
end
19'd1060: begin  
end
19'd1061: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd1062: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd1063: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd1064: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd1065: begin  
rid<=0;
end
19'd1201: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=7;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12447;
 end   
19'd1202: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=91;
   mapp<=50;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15127;
 end   
19'd1203: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=7;
   mapp<=41;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12633;
 end   
19'd1204: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=37;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd1205: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=57;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd1206: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=87;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd1207: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=53;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd1208: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=83;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd1209: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=22;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=21902;
 end   
19'd1210: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=46;
   mapp<=9;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=19703;
 end   
19'd1211: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=6;
   mapp<=9;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=25242;
 end   
19'd1212: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=30;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd1213: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=13;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd1214: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=68;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd1215: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd1216: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=91;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd1217: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd1359: begin  
rid<=1;
end
19'd1360: begin  
end
19'd1361: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd1362: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd1363: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd1364: begin  
rid<=0;
end
19'd1501: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=2;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11698;
 end   
19'd1502: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=50;
   mapp<=59;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=14465;
 end   
19'd1503: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=91;
   mapp<=24;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=17124;
 end   
19'd1504: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=36;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd1505: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=74;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd1506: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=20;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd1507: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd1508: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd1509: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=53;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=30883;
 end   
19'd1510: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=99;
   mapp<=21;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=31824;
 end   
19'd1511: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=18;
   mapp<=48;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=36877;
 end   
19'd1512: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=38;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd1513: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd1514: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=88;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd1515: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd1516: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd1517: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd1659: begin  
rid<=1;
end
19'd1660: begin  
end
19'd1661: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd1662: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd1663: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd1664: begin  
rid<=0;
end
19'd1801: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=16;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6893;
 end   
19'd1802: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=35;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8630;
 end   
19'd1803: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=51;
   mapp<=48;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4863;
 end   
19'd1804: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=83;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3754;
 end   
19'd1805: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=49;
   mapp<=7;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2300;
 end   
19'd1806: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=19;
   mapp<=21;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=2460;
 end   
19'd1807: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd1808: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd1809: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd1810: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd1811: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd1812: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=93;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=18716;
 end   
19'd1813: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=43;
   mapp<=98;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=19764;
 end   
19'd1814: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=23;
   mapp<=3;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=10579;
 end   
19'd1815: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=87;
   mapp<=24;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=9377;
 end   
19'd1816: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=14;
   mapp<=8;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=13199;
 end   
19'd1817: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=3;
   mapp<=44;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=10745;
 end   
19'd1818: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd1819: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd1820: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd1821: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd1822: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd1823: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd1965: begin  
rid<=1;
end
19'd1966: begin  
end
19'd1967: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd1968: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd1969: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd1970: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd1971: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd1972: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd1973: begin  
rid<=0;
end
19'd2101: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=80;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6368;
 end   
19'd2102: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=96;
   mapp<=18;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7342;
 end   
19'd2103: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=98;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7162;
 end   
19'd2104: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=81;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6330;
 end   
19'd2105: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=89;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6966;
 end   
19'd2106: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=98;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=5896;
 end   
19'd2107: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=9;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=1608;
 end   
19'd2108: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=57;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=4672;
 end   
19'd2109: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=72;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=4652;
 end   
19'd2110: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=22;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=2050;
 end   
19'd2111: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd2112: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=79;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17056;
 end   
19'd2113: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=90;
   mapp<=38;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=17788;
 end   
19'd2114: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=57;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=14610;
 end   
19'd2115: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=58;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=15124;
 end   
19'd2116: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=91;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=15908;
 end   
19'd2117: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=15;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=10620;
 end   
19'd2118: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=88;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=11832;
 end   
19'd2119: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=56;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=10242;
 end   
19'd2120: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=11;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=5740;
 end   
19'd2121: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=2;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=3526;
 end   
19'd2122: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd2123: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd2265: begin  
rid<=1;
end
19'd2266: begin  
end
19'd2267: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd2268: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd2269: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd2270: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd2271: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd2272: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd2273: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd2274: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd2275: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd2276: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd2277: begin  
rid<=0;
end
19'd2401: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=42;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4192;
 end   
19'd2402: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=44;
   mapp<=46;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6046;
 end   
19'd2403: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=16;
   mapp<=62;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7608;
 end   
19'd2404: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=86;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7470;
 end   
19'd2405: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=75;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5746;
 end   
19'd2406: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd2407: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd2408: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=76;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=21322;
 end   
19'd2409: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=92;
   mapp<=98;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20057;
 end   
19'd2410: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=89;
   mapp<=22;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15841;
 end   
19'd2411: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=51;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=22089;
 end   
19'd2412: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=21;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=21523;
 end   
19'd2413: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd2414: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd2415: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd2557: begin  
rid<=1;
end
19'd2558: begin  
end
19'd2559: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd2560: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd2561: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd2562: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd2563: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd2564: begin  
rid<=0;
end
19'd2701: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5475;
 end   
19'd2702: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=1;
   mapp<=10;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2774;
 end   
19'd2703: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=89;
   mapp<=3;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5962;
 end   
19'd2704: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=55;
   mapp<=69;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=11133;
 end   
19'd2705: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=23;
   mapp<=61;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=11158;
 end   
19'd2706: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=2;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=12379;
 end   
19'd2707: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=85;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd2708: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=82;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd2709: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=85;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd2710: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd2711: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=69;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14664;
 end   
19'd2712: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=54;
   mapp<=17;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12968;
 end   
19'd2713: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=21;
   mapp<=57;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15457;
 end   
19'd2714: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=89;
   mapp<=32;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=21512;
 end   
19'd2715: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=76;
   mapp<=32;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=21247;
 end   
19'd2716: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=29;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=22093;
 end   
19'd2717: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=68;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd2718: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=92;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd2719: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=25;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd2720: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=55;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd2721: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd2863: begin  
rid<=1;
end
19'd2864: begin  
end
19'd2865: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd2866: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd2867: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd2868: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd2869: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd2870: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd2871: begin  
rid<=0;
end
19'd3001: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=60;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5061;
 end   
19'd3002: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=18;
   mapp<=12;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3139;
 end   
19'd3003: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=53;
   mapp<=45;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3696;
 end   
19'd3004: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=39;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5460;
 end   
19'd3005: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd3006: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=79;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd3007: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=49;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14898;
 end   
19'd3008: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=37;
   mapp<=87;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=13854;
 end   
19'd3009: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=66;
   mapp<=29;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=16992;
 end   
19'd3010: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=49;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=21010;
 end   
19'd3011: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=93;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd3012: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=95;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd3013: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd3155: begin  
rid<=1;
end
19'd3156: begin  
end
19'd3157: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd3158: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd3159: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd3160: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd3161: begin  
rid<=0;
end
19'd3301: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=71;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6106;
 end   
19'd3302: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=365;
 end   
19'd3303: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=88;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6268;
 end   
19'd3304: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=82;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5852;
 end   
19'd3305: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=55;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3945;
 end   
19'd3306: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=34;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=2464;
 end   
19'd3307: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=14;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=1054;
 end   
19'd3308: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=1;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=141;
 end   
19'd3309: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=16;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=1216;
 end   
19'd3310: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=45;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=9976;
 end   
19'd3311: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=63;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=3200;
 end   
19'd3312: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=13;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=6853;
 end   
19'd3313: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=55;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=8327;
 end   
19'd3314: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=85;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=7770;
 end   
19'd3315: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=53;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=4849;
 end   
19'd3316: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=12;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=1594;
 end   
19'd3317: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=8;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=501;
 end   
19'd3318: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=32;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=2656;
 end   
19'd3319: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd3461: begin  
rid<=1;
end
19'd3462: begin  
end
19'd3463: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd3464: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd3465: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd3466: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd3467: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd3468: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd3469: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd3470: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd3471: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd3472: begin  
rid<=0;
end
19'd3601: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=46;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5722;
 end   
19'd3602: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=82;
   mapp<=58;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6430;
 end   
19'd3603: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=81;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4273;
 end   
19'd3604: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=44;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd3605: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=29;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=9848;
 end   
19'd3606: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=61;
   mapp<=22;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=13056;
 end   
19'd3607: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=35;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=8733;
 end   
19'd3608: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=50;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd3609: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd3751: begin  
rid<=1;
end
19'd3752: begin  
end
19'd3753: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd3754: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd3755: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd3756: begin  
rid<=0;
end
19'd3901: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=49;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14110;
 end   
19'd3902: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=86;
   mapp<=59;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=19442;
 end   
19'd3903: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=13;
   mapp<=92;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12215;
 end   
19'd3904: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=74;
   mapp<=39;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=14087;
 end   
19'd3905: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=22;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd3906: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=68;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd3907: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd3908: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd3909: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd3910: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=14;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=27582;
 end   
19'd3911: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=24;
   mapp<=87;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=31105;
 end   
19'd3912: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=34;
   mapp<=5;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=23262;
 end   
19'd3913: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=74;
   mapp<=58;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=25371;
 end   
19'd3914: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=72;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd3915: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=59;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd3916: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd3917: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd3918: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd3919: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd4061: begin  
rid<=1;
end
19'd4062: begin  
end
19'd4063: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd4064: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd4065: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd4066: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd4067: begin  
rid<=0;
end
19'd4201: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=85;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=22514;
 end   
19'd4202: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=2;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=24690;
 end   
19'd4203: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=80;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd4204: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=13;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd4205: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=27;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd4206: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=2;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd4207: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=99;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd4208: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=27;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd4209: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=25;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd4210: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=43;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd4211: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=25;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=45192;
 end   
19'd4212: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=31;
   mapp<=23;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=45089;
 end   
19'd4213: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=92;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd4214: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=42;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd4215: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=22;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd4216: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=86;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd4217: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=64;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd4218: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd4219: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=87;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd4220: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=60;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd4221: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd4363: begin  
rid<=1;
end
19'd4364: begin  
end
19'd4365: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd4366: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd4367: begin  
rid<=0;
end
19'd4501: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=67;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=22748;
 end   
19'd4502: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=85;
   mapp<=70;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=18271;
 end   
19'd4503: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=50;
   mapp<=35;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=16549;
 end   
19'd4504: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=40;
   mapp<=33;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=22532;
 end   
19'd4505: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=94;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd4506: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=95;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd4507: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=24;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd4508: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=19;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd4509: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=25;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd4510: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=76;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd4511: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=51;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=42304;
 end   
19'd4512: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=84;
   mapp<=58;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=40211;
 end   
19'd4513: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=18;
   mapp<=2;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=38049;
 end   
19'd4514: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=64;
   mapp<=71;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=42594;
 end   
19'd4515: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=19;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd4516: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=52;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd4517: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd4518: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=87;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd4519: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=60;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd4520: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=26;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd4521: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd4663: begin  
rid<=1;
end
19'd4664: begin  
end
19'd4665: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd4666: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd4667: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd4668: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd4669: begin  
rid<=0;
end
19'd4801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=76;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5725;
 end   
19'd4802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=27;
   mapp<=15;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2545;
 end   
19'd4803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=43;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3900;
 end   
19'd4804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=58;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5050;
 end   
19'd4805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=64;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4655;
 end   
19'd4806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=9;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd4807: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=65;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=18537;
 end   
19'd4808: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=87;
   mapp<=86;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=16301;
 end   
19'd4809: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=77;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=16578;
 end   
19'd4810: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=74;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=13268;
 end   
19'd4811: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=25;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=9027;
 end   
19'd4812: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=27;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd4813: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd4955: begin  
rid<=1;
end
19'd4956: begin  
end
19'd4957: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd4958: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd4959: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd4960: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd4961: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd4962: begin  
rid<=0;
end
19'd5101: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=25;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6309;
 end   
19'd5102: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=64;
   mapp<=20;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8636;
 end   
19'd5103: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=60;
   mapp<=2;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10502;
 end   
19'd5104: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=2;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd5105: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=16;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd5106: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=30;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd5107: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=26;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd5108: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd5109: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd5110: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=63;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16024;
 end   
19'd5111: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=40;
   mapp<=71;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20124;
 end   
19'd5112: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=51;
   mapp<=11;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=20772;
 end   
19'd5113: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=62;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd5114: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=29;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd5115: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd5116: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=13;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd5117: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd5118: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd5119: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd5261: begin  
rid<=1;
end
19'd5262: begin  
end
19'd5263: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd5264: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd5265: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd5266: begin  
rid<=0;
end
19'd5401: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=3;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=195;
 end   
19'd5402: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=7;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=31;
 end   
19'd5403: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=77;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=251;
 end   
19'd5404: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=30;
 end   
19'd5405: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=58;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=214;
 end   
19'd5406: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=39;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=167;
 end   
19'd5407: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=87;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5415;
 end   
19'd5408: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=57;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=4990;
 end   
19'd5409: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=24;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=2339;
 end   
19'd5410: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=77;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6729;
 end   
19'd5411: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=8;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=910;
 end   
19'd5412: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=13;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=1298;
 end   
19'd5413: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd5555: begin  
rid<=1;
end
19'd5556: begin  
end
19'd5557: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd5558: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd5559: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd5560: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd5561: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd5562: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd5563: begin  
rid<=0;
end
19'd5701: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=93;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7932;
 end   
19'd5702: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=84;
   mapp<=28;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5190;
 end   
19'd5703: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=5;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1440;
 end   
19'd5704: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=40;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd5705: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=35;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8541;
 end   
19'd5706: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=56;
   mapp<=4;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=6094;
 end   
19'd5707: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=72;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=2432;
 end   
19'd5708: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=50;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd5709: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd5851: begin  
rid<=1;
end
19'd5852: begin  
end
19'd5853: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd5854: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd5855: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd5856: begin  
rid<=0;
end
19'd6001: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=57;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5090;
 end   
19'd6002: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=26;
   mapp<=16;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3340;
 end   
19'd6003: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=57;
   mapp<=26;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5650;
 end   
19'd6004: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=37;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5032;
 end   
19'd6005: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=71;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6706;
 end   
19'd6006: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=69;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7386;
 end   
19'd6007: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=61;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=5584;
 end   
19'd6008: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=96;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=6240;
 end   
19'd6009: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=22;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd6010: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=17;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd6011: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=85;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=9015;
 end   
19'd6012: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=41;
   mapp<=17;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=7007;
 end   
19'd6013: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=23;
   mapp<=96;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=9203;
 end   
19'd6014: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=29;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=12113;
 end   
19'd6015: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=29;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=13823;
 end   
19'd6016: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=65;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=12241;
 end   
19'd6017: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=59;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=16052;
 end   
19'd6018: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=32;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=13536;
 end   
19'd6019: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=96;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd6020: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=55;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd6021: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd6163: begin  
rid<=1;
end
19'd6164: begin  
end
19'd6165: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd6166: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd6167: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd6168: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd6169: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd6170: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd6171: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd6172: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd6173: begin  
rid<=0;
end
19'd6301: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=83;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6972;
 end   
19'd6302: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=34;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2832;
 end   
19'd6303: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=54;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4502;
 end   
19'd6304: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=72;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6006;
 end   
19'd6305: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=57;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4771;
 end   
19'd6306: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=69;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=5777;
 end   
19'd6307: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=32;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=2716;
 end   
19'd6308: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=63;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=5299;
 end   
19'd6309: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=7;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=661;
 end   
19'd6310: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=11;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7093;
 end   
19'd6311: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=3217;
 end   
19'd6312: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=67;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=5239;
 end   
19'd6313: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=48;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6534;
 end   
19'd6314: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=75;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=5596;
 end   
19'd6315: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=38;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=6195;
 end   
19'd6316: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=23;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=2969;
 end   
19'd6317: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=42;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=5761;
 end   
19'd6318: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=54;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=1255;
 end   
19'd6319: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd6461: begin  
rid<=1;
end
19'd6462: begin  
end
19'd6463: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd6464: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd6465: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd6466: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd6467: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd6468: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd6469: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd6470: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd6471: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd6472: begin  
rid<=0;
end
19'd6601: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=34;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2131;
 end   
19'd6602: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=5;
   mapp<=25;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=965;
 end   
19'd6603: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=21;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1084;
 end   
19'd6604: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=70;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=2540;
 end   
19'd6605: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd6606: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=93;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=11550;
 end   
19'd6607: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=34;
   mapp<=50;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8947;
 end   
19'd6608: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=98;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=12884;
 end   
19'd6609: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=79;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=9921;
 end   
19'd6610: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd6611: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd6753: begin  
rid<=1;
end
19'd6754: begin  
end
19'd6755: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd6756: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd6757: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd6758: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd6759: begin  
rid<=0;
end
19'd6901: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=55;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11387;
 end   
19'd6902: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=55;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9515;
 end   
19'd6903: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=42;
   mapp<=76;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7079;
 end   
19'd6904: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=5;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5731;
 end   
19'd6905: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=62;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=9492;
 end   
19'd6906: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=48;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7145;
 end   
19'd6907: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=81;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=5061;
 end   
19'd6908: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=2507;
 end   
19'd6909: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd6910: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd6911: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=13;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=18562;
 end   
19'd6912: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=75;
   mapp<=11;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=17161;
 end   
19'd6913: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=72;
   mapp<=77;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15496;
 end   
19'd6914: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=24;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=15637;
 end   
19'd6915: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=78;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=17502;
 end   
19'd6916: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=52;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=17958;
 end   
19'd6917: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=43;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=18076;
 end   
19'd6918: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=96;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=12110;
 end   
19'd6919: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd6920: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd6921: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd7063: begin  
rid<=1;
end
19'd7064: begin  
end
19'd7065: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd7066: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd7067: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd7068: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd7069: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd7070: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd7071: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd7072: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd7073: begin  
rid<=0;
end
19'd7201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=69;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11005;
 end   
19'd7202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=31;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10948;
 end   
19'd7203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=40;
   mapp<=12;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=13086;
 end   
19'd7204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=88;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd7205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=85;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd7206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=90;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd7207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=53;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=23782;
 end   
19'd7208: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=14;
   mapp<=89;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=22425;
 end   
19'd7209: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=51;
   mapp<=90;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=28163;
 end   
19'd7210: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=40;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd7211: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=44;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd7212: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=58;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd7213: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd7355: begin  
rid<=1;
end
19'd7356: begin  
end
19'd7357: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd7358: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd7359: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd7360: begin  
rid<=0;
end
19'd7501: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=75;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=20685;
 end   
19'd7502: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=8;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8640;
 end   
19'd7503: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=92;
   mapp<=64;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8557;
 end   
19'd7504: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=97;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd7505: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd7506: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd7507: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=29;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=27137;
 end   
19'd7508: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=40;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18013;
 end   
19'd7509: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=13;
   mapp<=61;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15311;
 end   
19'd7510: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=74;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd7511: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd7512: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd7513: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd7655: begin  
rid<=1;
end
19'd7656: begin  
end
19'd7657: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd7658: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd7659: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd7660: begin  
rid<=0;
end
19'd7801: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=27;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=18686;
 end   
19'd7802: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=84;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=18845;
 end   
19'd7803: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=75;
   mapp<=13;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=23131;
 end   
19'd7804: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=86;
   mapp<=92;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=23199;
 end   
19'd7805: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=98;
   mapp<=24;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=21566;
 end   
19'd7806: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=70;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd7807: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd7808: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd7809: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd7810: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd7811: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=89;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=29909;
 end   
19'd7812: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=40;
   mapp<=47;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=25537;
 end   
19'd7813: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=64;
   mapp<=4;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=28530;
 end   
19'd7814: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=42;
   mapp<=3;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=29917;
 end   
19'd7815: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=19;
   mapp<=21;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=30098;
 end   
19'd7816: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=13;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd7817: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd7818: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd7819: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd7820: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd7821: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd7963: begin  
rid<=1;
end
19'd7964: begin  
end
19'd7965: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd7966: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd7967: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd7968: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd7969: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd7970: begin  
rid<=0;
end
19'd8101: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=50;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1060;
 end   
19'd8102: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=5;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2500;
 end   
19'd8103: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=75;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2618;
 end   
19'd8104: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=39;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=828;
 end   
19'd8105: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=3;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=798;
 end   
19'd8106: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=22;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd8107: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=84;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=11548;
 end   
19'd8108: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=48;
   mapp<=47;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=10541;
 end   
19'd8109: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=71;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=12584;
 end   
19'd8110: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=64;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=7711;
 end   
19'd8111: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=13;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=5597;
 end   
19'd8112: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=75;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd8113: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd8255: begin  
rid<=1;
end
19'd8256: begin  
end
19'd8257: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd8258: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd8259: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd8260: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd8261: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd8262: begin  
rid<=0;
end
19'd8401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=65;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9215;
 end   
19'd8402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=40;
   mapp<=78;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10630;
 end   
19'd8403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=45;
   mapp<=69;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7840;
 end   
19'd8404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=62;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=8645;
 end   
19'd8405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=19;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=8680;
 end   
19'd8406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=85;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=11115;
 end   
19'd8407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd8408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd8409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=87;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=15581;
 end   
19'd8410: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=70;
   mapp<=18;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=17159;
 end   
19'd8411: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=63;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15449;
 end   
19'd8412: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=1;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=12358;
 end   
19'd8413: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=23;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=17457;
 end   
19'd8414: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=32;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=22215;
 end   
19'd8415: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd8416: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd8417: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd8559: begin  
rid<=1;
end
19'd8560: begin  
end
19'd8561: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd8562: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd8563: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd8564: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd8565: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd8566: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd8567: begin  
rid<=0;
end
19'd8701: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=15;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5067;
 end   
19'd8702: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=65;
   mapp<=27;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5504;
 end   
19'd8703: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=28;
   mapp<=0;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7897;
 end   
19'd8704: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=43;
   mapp<=69;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5255;
 end   
19'd8705: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=47;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6050;
 end   
19'd8706: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=88;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=3856;
 end   
19'd8707: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=43;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=6395;
 end   
19'd8708: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd8709: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=9;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd8710: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=63;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd8711: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=8;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14603;
 end   
19'd8712: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=60;
   mapp<=81;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=17517;
 end   
19'd8713: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=21;
   mapp<=88;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=22072;
 end   
19'd8714: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=58;
   mapp<=42;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=22147;
 end   
19'd8715: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=54;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=23652;
 end   
19'd8716: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=88;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=21872;
 end   
19'd8717: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=46;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=22057;
 end   
19'd8718: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=90;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd8719: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=49;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd8720: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=43;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd8721: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd8863: begin  
rid<=1;
end
19'd8864: begin  
end
19'd8865: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd8866: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd8867: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd8868: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd8869: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd8870: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd8871: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd8872: begin  
rid<=0;
end
19'd9001: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=83;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6329;
 end   
19'd9002: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=35;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6831;
 end   
19'd9003: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd9004: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=53;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=10172;
 end   
19'd9005: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=29;
   mapp<=85;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12438;
 end   
19'd9006: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd9007: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd9149: begin  
rid<=1;
end
19'd9150: begin  
end
19'd9151: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd9152: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd9153: begin  
rid<=0;
end
19'd9301: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=55;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5635;
 end   
19'd9302: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=18;
   mapp<=59;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6655;
 end   
19'd9303: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=26;
   mapp<=57;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6366;
 end   
19'd9304: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=11;
   mapp<=66;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7115;
 end   
19'd9305: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=25;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd9306: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=55;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd9307: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=1;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd9308: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=49;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd9309: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=75;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=22717;
 end   
19'd9310: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=13;
   mapp<=84;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18967;
 end   
19'd9311: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=42;
   mapp<=15;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=24882;
 end   
19'd9312: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=96;
   mapp<=64;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=23359;
 end   
19'd9313: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=48;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd9314: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=72;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd9315: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=26;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd9316: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=6;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd9317: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd9459: begin  
rid<=1;
end
19'd9460: begin  
end
19'd9461: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd9462: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd9463: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd9464: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd9465: begin  
rid<=0;
end
19'd9601: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=93;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5140;
 end   
19'd9602: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=65;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2928;
 end   
19'd9603: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=36;
   mapp<=26;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8628;
 end   
19'd9604: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=36;
   mapp<=12;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6071;
 end   
19'd9605: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=41;
   mapp<=75;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=7290;
 end   
19'd9606: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=14;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=5356;
 end   
19'd9607: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=94;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd9608: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=56;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd9609: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=52;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd9610: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=36;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd9611: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=30;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12329;
 end   
19'd9612: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=41;
   mapp<=82;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=10362;
 end   
19'd9613: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=25;
   mapp<=55;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=16595;
 end   
19'd9614: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=11;
   mapp<=15;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=17153;
 end   
19'd9615: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=37;
   mapp<=31;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=23370;
 end   
19'd9616: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=86;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=20738;
 end   
19'd9617: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=90;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd9618: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=50;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd9619: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd9620: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd9621: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd9763: begin  
rid<=1;
end
19'd9764: begin  
end
19'd9765: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd9766: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd9767: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd9768: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd9769: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd9770: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd9771: begin  
rid<=0;
end
19'd9901: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=33;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3360;
 end   
19'd9902: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=54;
   mapp<=52;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2344;
 end   
19'd9903: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=3;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd9904: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd9905: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=24;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=4955;
 end   
19'd9906: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=17;
   mapp<=3;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=3992;
 end   
19'd9907: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=13;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd9908: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd9909: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd10051: begin  
rid<=1;
end
19'd10052: begin  
end
19'd10053: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd10054: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd10055: begin  
rid<=0;
end
19'd10201: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=61;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11732;
 end   
19'd10202: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=64;
   mapp<=80;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12381;
 end   
19'd10203: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=3;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd10204: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=76;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd10205: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=43;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd10206: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd10207: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=53;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14859;
 end   
19'd10208: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=74;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20763;
 end   
19'd10209: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=20;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd10210: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=2;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd10211: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=23;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd10212: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd10213: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd10355: begin  
rid<=1;
end
19'd10356: begin  
end
19'd10357: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd10358: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd10359: begin  
rid<=0;
end
19'd10501: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=71;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7614;
 end   
19'd10502: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=3;
   mapp<=59;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3623;
 end   
19'd10503: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=45;
   mapp<=8;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10089;
 end   
19'd10504: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=81;
   mapp<=19;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=8935;
 end   
19'd10505: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=4;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6707;
 end   
19'd10506: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=92;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=14207;
 end   
19'd10507: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=85;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=9932;
 end   
19'd10508: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=13;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd10509: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=98;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd10510: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd10511: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=61;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=11154;
 end   
19'd10512: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=34;
   mapp<=38;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=7522;
 end   
19'd10513: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=8;
   mapp<=37;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15696;
 end   
19'd10514: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=61;
   mapp<=10;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=16110;
 end   
19'd10515: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=59;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=12784;
 end   
19'd10516: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=93;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=19746;
 end   
19'd10517: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=15;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=14943;
 end   
19'd10518: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=69;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd10519: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd10520: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=69;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd10521: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd10663: begin  
rid<=1;
end
19'd10664: begin  
end
19'd10665: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd10666: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd10667: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd10668: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd10669: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd10670: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd10671: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd10672: begin  
rid<=0;
end
19'd10801: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=55;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5960;
 end   
19'd10802: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=15;
   mapp<=64;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3838;
 end   
19'd10803: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=30;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd10804: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=39;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd10805: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd10806: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=10;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=24524;
 end   
19'd10807: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=84;
   mapp<=82;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=22893;
 end   
19'd10808: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=74;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd10809: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=80;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd10810: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=15;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd10811: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd10953: begin  
rid<=1;
end
19'd10954: begin  
end
19'd10955: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd10956: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd10957: begin  
rid<=0;
end
19'd11101: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=98;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8117;
 end   
19'd11102: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=73;
   mapp<=79;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8827;
 end   
19'd11103: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=88;
   mapp<=10;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7743;
 end   
19'd11104: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=77;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4273;
 end   
19'd11105: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=32;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5834;
 end   
19'd11106: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=56;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=8051;
 end   
19'd11107: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd11108: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=13;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd11109: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=23;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=13404;
 end   
19'd11110: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=63;
   mapp<=41;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18039;
 end   
19'd11111: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=28;
   mapp<=90;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=18431;
 end   
19'd11112: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=84;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=8143;
 end   
19'd11113: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=78;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=12848;
 end   
19'd11114: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=18612;
 end   
19'd11115: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=71;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd11116: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=85;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd11117: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd11259: begin  
rid<=1;
end
19'd11260: begin  
end
19'd11261: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd11262: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd11263: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd11264: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd11265: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd11266: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd11267: begin  
rid<=0;
end
19'd11401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=50;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=23376;
 end   
19'd11402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=98;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=17883;
 end   
19'd11403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=9;
   mapp<=53;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=21453;
 end   
19'd11404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=93;
   mapp<=95;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=21231;
 end   
19'd11405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=86;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd11406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd11407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd11408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd11409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=5;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=26776;
 end   
19'd11410: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=26;
   mapp<=16;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=22811;
 end   
19'd11411: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=16;
   mapp<=49;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=26816;
 end   
19'd11412: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=16;
   mapp<=67;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=25128;
 end   
19'd11413: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=26;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd11414: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd11415: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd11416: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd11417: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd11559: begin  
rid<=1;
end
19'd11560: begin  
end
19'd11561: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd11562: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd11563: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd11564: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd11565: begin  
rid<=0;
end
19'd11701: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=64;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5184;
 end   
19'd11702: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=40;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3250;
 end   
19'd11703: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=86;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6986;
 end   
19'd11704: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=21;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1731;
 end   
19'd11705: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=21;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=6486;
 end   
19'd11706: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=64;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=7218;
 end   
19'd11707: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=9;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=7544;
 end   
19'd11708: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=15;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=2661;
 end   
19'd11709: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd11851: begin  
rid<=1;
end
19'd11852: begin  
end
19'd11853: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd11854: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd11855: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd11856: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd11857: begin  
rid<=0;
end
19'd12001: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=6;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4244;
 end   
19'd12002: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=68;
   mapp<=41;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5576;
 end   
19'd12003: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=18;
   mapp<=45;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3518;
 end   
19'd12004: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=2;
   mapp<=62;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7094;
 end   
19'd12005: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=7;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd12006: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=7;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd12007: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=81;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd12008: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd12009: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=36;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd12010: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=93;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16622;
 end   
19'd12011: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=96;
   mapp<=14;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18218;
 end   
19'd12012: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=52;
   mapp<=9;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=17789;
 end   
19'd12013: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=54;
   mapp<=84;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=19624;
 end   
19'd12014: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=45;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd12015: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=8;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd12016: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=48;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd12017: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=91;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd12018: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd12019: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd12161: begin  
rid<=1;
end
19'd12162: begin  
end
19'd12163: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd12164: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd12165: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd12166: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd12167: begin  
rid<=0;
end
19'd12301: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=69;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13343;
 end   
19'd12302: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=79;
   mapp<=58;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15211;
 end   
19'd12303: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=38;
   mapp<=22;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=14197;
 end   
19'd12304: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=23;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd12305: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=18;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd12306: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=66;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd12307: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=59;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd12308: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=98;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd12309: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=46;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=33252;
 end   
19'd12310: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=92;
   mapp<=96;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=33184;
 end   
19'd12311: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=37;
   mapp<=62;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=24877;
 end   
19'd12312: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=25;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd12313: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=47;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd12314: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=58;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd12315: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=2;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd12316: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=7;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd12317: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd12459: begin  
rid<=1;
end
19'd12460: begin  
end
19'd12461: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd12462: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd12463: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd12464: begin  
rid<=0;
end
19'd12601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=40;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3680;
 end   
19'd12602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10;
 end   
19'd12603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=78;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3140;
 end   
19'd12604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=99;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3990;
 end   
19'd12605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=52;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2120;
 end   
19'd12606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=48;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=1970;
 end   
19'd12607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=82;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=3340;
 end   
19'd12608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=97;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5135;
 end   
19'd12609: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=75;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=7285;
 end   
19'd12610: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=62;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=9154;
 end   
19'd12611: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=67;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=10489;
 end   
19'd12612: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=36;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=5612;
 end   
19'd12613: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=97;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=11379;
 end   
19'd12614: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=18;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=5086;
 end   
19'd12615: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd12757: begin  
rid<=1;
end
19'd12758: begin  
end
19'd12759: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd12760: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd12761: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd12762: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd12763: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd12764: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd12765: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd12766: begin  
rid<=0;
end
19'd12901: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=30;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=480;
 end   
19'd12902: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=49;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=794;
 end   
19'd12903: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=25;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=420;
 end   
19'd12904: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=29;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=2162;
 end   
19'd12905: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=20;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=1954;
 end   
19'd12906: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=40;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=2740;
 end   
19'd12907: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd13049: begin  
rid<=1;
end
19'd13050: begin  
end
19'd13051: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd13052: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd13053: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd13054: begin  
rid<=0;
end
19'd13201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=61;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3782;
 end   
19'd13202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=55;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3365;
 end   
19'd13203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=75;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4595;
 end   
19'd13204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=92;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5642;
 end   
19'd13205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=46;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=6266;
 end   
19'd13206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=98;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=7873;
 end   
19'd13207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=46;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=6711;
 end   
19'd13208: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=14;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6286;
 end   
19'd13209: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd13351: begin  
rid<=1;
end
19'd13352: begin  
end
19'd13353: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd13354: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd13355: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd13356: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd13357: begin  
rid<=0;
end
19'd13501: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=15;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=570;
 end   
19'd13502: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=63;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=955;
 end   
19'd13503: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=75;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1145;
 end   
19'd13504: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=28;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=1158;
 end   
19'd13505: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=75;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=3055;
 end   
19'd13506: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=15;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=1565;
 end   
19'd13507: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd13649: begin  
rid<=1;
end
19'd13650: begin  
end
19'd13651: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd13652: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd13653: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd13654: begin  
rid<=0;
end
19'd13801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=57;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4253;
 end   
19'd13802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=62;
   mapp<=64;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4224;
 end   
19'd13803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=61;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1861;
 end   
19'd13804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=24;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3286;
 end   
19'd13805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=49;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4701;
 end   
19'd13806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=69;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=2315;
 end   
19'd13807: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=30;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=1682;
 end   
19'd13808: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=23;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=3385;
 end   
19'd13809: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=50;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd13810: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=10;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5508;
 end   
19'd13811: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=37;
   mapp<=25;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=6345;
 end   
19'd13812: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=36;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=3974;
 end   
19'd13813: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=37;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6457;
 end   
19'd13814: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=78;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=9600;
 end   
19'd13815: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=93;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=6284;
 end   
19'd13816: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=36;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=3220;
 end   
19'd13817: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=14;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=5447;
 end   
19'd13818: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=64;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd13819: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd13961: begin  
rid<=1;
end
19'd13962: begin  
end
19'd13963: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd13964: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd13965: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd13966: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd13967: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd13968: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd13969: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd13970: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd13971: begin  
rid<=0;
end
19'd14101: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=85;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13034;
 end   
19'd14102: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=52;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=13421;
 end   
19'd14103: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=73;
   mapp<=37;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=18814;
 end   
19'd14104: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=52;
   mapp<=4;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=16257;
 end   
19'd14105: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=94;
   mapp<=37;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=20719;
 end   
19'd14106: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=76;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd14107: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=26;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd14108: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd14109: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd14110: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd14111: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd14112: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=65;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=28811;
 end   
19'd14113: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=5;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=24624;
 end   
19'd14114: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=85;
   mapp<=49;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=31477;
 end   
19'd14115: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=16;
   mapp<=40;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=23496;
 end   
19'd14116: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=50;
   mapp<=74;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=33011;
 end   
19'd14117: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=15;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd14118: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=9;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd14119: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd14120: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd14121: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd14122: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd14123: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd14265: begin  
rid<=1;
end
19'd14266: begin  
end
19'd14267: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd14268: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd14269: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd14270: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd14271: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd14272: begin  
rid<=0;
end
19'd14401: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=58;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8300;
 end   
19'd14402: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=31;
   mapp<=74;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7051;
 end   
19'd14403: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=68;
   mapp<=9;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8900;
 end   
19'd14404: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=26;
   mapp<=0;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=10253;
 end   
19'd14405: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=95;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=15451;
 end   
19'd14406: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=73;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=13063;
 end   
19'd14407: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=89;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=13777;
 end   
19'd14408: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd14409: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd14410: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd14411: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=74;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14941;
 end   
19'd14412: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=64;
   mapp<=22;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=14123;
 end   
19'd14413: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=2;
   mapp<=74;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=22312;
 end   
19'd14414: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=55;
   mapp<=79;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=21353;
 end   
19'd14415: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=10;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=24688;
 end   
19'd14416: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=52;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=27566;
 end   
19'd14417: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=82;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=29379;
 end   
19'd14418: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd14419: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd14420: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd14421: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd14563: begin  
rid<=1;
end
19'd14564: begin  
end
19'd14565: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd14566: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd14567: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd14568: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd14569: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd14570: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd14571: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd14572: begin  
rid<=0;
end
19'd14701: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=5;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2355;
 end   
19'd14702: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=95;
   mapp<=21;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2205;
 end   
19'd14703: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=22;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4595;
 end   
19'd14704: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=47;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7580;
 end   
19'd14705: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=77;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=8880;
 end   
19'd14706: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd14707: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=72;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=11073;
 end   
19'd14708: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=39;
   mapp<=50;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=7482;
 end   
19'd14709: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=43;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=9797;
 end   
19'd14710: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=54;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=14627;
 end   
19'd14711: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=81;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=15180;
 end   
19'd14712: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd14713: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd14855: begin  
rid<=1;
end
19'd14856: begin  
end
19'd14857: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd14858: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd14859: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd14860: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd14861: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd14862: begin  
rid<=0;
end
19'd15001: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=86;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9310;
 end   
19'd15002: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=19;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11186;
 end   
19'd15003: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=58;
   mapp<=8;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5090;
 end   
19'd15004: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=45;
   mapp<=15;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5929;
 end   
19'd15005: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=6;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd15006: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=66;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd15007: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd15008: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd15009: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd15010: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=83;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=25592;
 end   
19'd15011: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=22;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=32100;
 end   
19'd15012: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=31;
   mapp<=92;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=28286;
 end   
19'd15013: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=76;
   mapp<=87;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=26123;
 end   
19'd15014: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=83;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd15015: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=48;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd15016: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd15017: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd15018: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd15019: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd15161: begin  
rid<=1;
end
19'd15162: begin  
end
19'd15163: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd15164: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd15165: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd15166: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd15167: begin  
rid<=0;
end
19'd15301: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=24;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=23327;
 end   
19'd15302: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=86;
   mapp<=76;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=24183;
 end   
19'd15303: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=77;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd15304: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=69;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd15305: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=43;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd15306: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=34;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd15307: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=77;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd15308: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=68;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd15309: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=68;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd15310: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=12;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=38316;
 end   
19'd15311: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=3;
   mapp<=96;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=37685;
 end   
19'd15312: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=27;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd15313: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=8;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd15314: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=45;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd15315: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=8;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd15316: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=85;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd15317: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=38;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd15318: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd15319: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd15461: begin  
rid<=1;
end
19'd15462: begin  
end
19'd15463: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd15464: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd15465: begin  
rid<=0;
end
19'd15601: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=67;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13583;
 end   
19'd15602: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=13;
   mapp<=50;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=18219;
 end   
19'd15603: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=93;
   mapp<=28;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=20937;
 end   
19'd15604: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=34;
   mapp<=11;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=20388;
 end   
19'd15605: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=72;
   mapp<=50;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=27169;
 end   
19'd15606: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=72;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd15607: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=30;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd15608: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd15609: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd15610: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd15611: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd15612: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=23;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=32166;
 end   
19'd15613: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=79;
   mapp<=42;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=40965;
 end   
19'd15614: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=95;
   mapp<=77;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=41609;
 end   
19'd15615: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=69;
   mapp<=77;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=38492;
 end   
19'd15616: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=27;
   mapp<=70;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=44372;
 end   
19'd15617: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=42;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd15618: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=10;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd15619: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd15620: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd15621: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd15622: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd15623: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd15765: begin  
rid<=1;
end
19'd15766: begin  
end
19'd15767: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd15768: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd15769: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd15770: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd15771: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd15772: begin  
rid<=0;
end
19'd15901: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=87;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2262;
 end   
19'd15902: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=70;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1830;
 end   
19'd15903: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=28;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=748;
 end   
19'd15904: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=51;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1356;
 end   
19'd15905: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=13;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=3016;
 end   
19'd15906: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=60;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=5310;
 end   
19'd15907: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=83;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=5562;
 end   
19'd15908: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=86;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6344;
 end   
19'd15909: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd16051: begin  
rid<=1;
end
19'd16052: begin  
end
19'd16053: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd16054: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd16055: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd16056: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd16057: begin  
rid<=0;
end
19'd16201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=18;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6323;
 end   
19'd16202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=3;
   mapp<=28;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5870;
 end   
19'd16203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=67;
   mapp<=34;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11277;
 end   
19'd16204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=65;
   mapp<=41;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=10865;
 end   
19'd16205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=38;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=9032;
 end   
19'd16206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=81;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=9752;
 end   
19'd16207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=57;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd16208: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=50;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd16209: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=14;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd16210: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=56;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=22582;
 end   
19'd16211: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=7;
   mapp<=58;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18714;
 end   
19'd16212: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=78;
   mapp<=61;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=30313;
 end   
19'd16213: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=89;
   mapp<=63;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=30307;
 end   
19'd16214: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=35;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=26225;
 end   
19'd16215: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=65;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=31136;
 end   
19'd16216: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=75;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd16217: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=86;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd16218: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=86;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd16219: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd16361: begin  
rid<=1;
end
19'd16362: begin  
end
19'd16363: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd16364: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd16365: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd16366: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd16367: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd16368: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd16369: begin  
rid<=0;
end
19'd16501: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=28;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=840;
 end   
19'd16502: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=0;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1354;
 end   
19'd16503: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=40;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=4520;
 end   
19'd16504: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=0;
   mapp<=33;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=2674;
 end   
19'd16505: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd16647: begin  
rid<=1;
end
19'd16648: begin  
end
19'd16649: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd16650: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd16651: begin  
rid<=0;
end
19'd16801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=37;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9478;
 end   
19'd16802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=92;
   mapp<=99;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9048;
 end   
19'd16803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=82;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3612;
 end   
19'd16804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=28;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5458;
 end   
19'd16805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=52;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=7391;
 end   
19'd16806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=69;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=5096;
 end   
19'd16807: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=44;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=9806;
 end   
19'd16808: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=94;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=1802;
 end   
19'd16809: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=8;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd16810: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=32;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12787;
 end   
19'd16811: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=35;
   mapp<=47;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=11244;
 end   
19'd16812: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=8;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=7036;
 end   
19'd16813: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=64;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=13345;
 end   
19'd16814: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=97;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=14456;
 end   
19'd16815: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=43;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=9635;
 end   
19'd16816: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=49;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=13059;
 end   
19'd16817: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=15;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=4509;
 end   
19'd16818: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=41;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd16819: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd16961: begin  
rid<=1;
end
19'd16962: begin  
end
19'd16963: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd16964: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd16965: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd16966: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd16967: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd16968: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd16969: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd16970: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd16971: begin  
rid<=0;
end
19'd17101: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=51;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4923;
 end   
19'd17102: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=74;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4575;
 end   
19'd17103: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=33;
   mapp<=23;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4784;
 end   
19'd17104: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=91;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=2364;
 end   
19'd17105: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4702;
 end   
19'd17106: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=54;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7249;
 end   
19'd17107: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=90;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd17108: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=97;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd17109: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=31;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12152;
 end   
19'd17110: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=44;
   mapp<=80;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=15397;
 end   
19'd17111: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=40;
   mapp<=78;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=20226;
 end   
19'd17112: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=87;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=13887;
 end   
19'd17113: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=99;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=15057;
 end   
19'd17114: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=25;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=17328;
 end   
19'd17115: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=83;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd17116: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd17117: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd17259: begin  
rid<=1;
end
19'd17260: begin  
end
19'd17261: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd17262: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd17263: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd17264: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd17265: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd17266: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd17267: begin  
rid<=0;
end
19'd17401: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=60;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3120;
 end   
19'd17402: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=0;
   mapp<=11;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=670;
 end   
19'd17403: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=97;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=6418;
 end   
19'd17404: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=0;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=4550;
 end   
19'd17405: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd17547: begin  
rid<=1;
end
19'd17548: begin  
end
19'd17549: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd17550: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd17551: begin  
rid<=0;
end
19'd17701: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=92;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8189;
 end   
19'd17702: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=10;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7753;
 end   
19'd17703: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=49;
   mapp<=91;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9559;
 end   
19'd17704: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=78;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=10006;
 end   
19'd17705: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=79;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd17706: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=71;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd17707: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=20;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=19228;
 end   
19'd17708: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=97;
   mapp<=73;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=24188;
 end   
19'd17709: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=26;
   mapp<=93;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=25479;
 end   
19'd17710: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=76;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=30054;
 end   
19'd17711: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=90;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd17712: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=82;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd17713: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd17855: begin  
rid<=1;
end
19'd17856: begin  
end
19'd17857: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd17858: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd17859: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd17860: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd17861: begin  
rid<=0;
end
19'd18001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=72;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12363;
 end   
19'd18002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=80;
   mapp<=89;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8355;
 end   
19'd18003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=8;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd18004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=67;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd18005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=8;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd18006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=77;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd18007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=22;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=23332;
 end   
19'd18008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=11;
   mapp<=70;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=22181;
 end   
19'd18009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=19;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd18010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=61;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd18011: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=56;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd18012: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=90;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd18013: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd18155: begin  
rid<=1;
end
19'd18156: begin  
end
19'd18157: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd18158: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd18159: begin  
rid<=0;
end
19'd18301: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=32;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=512;
 end   
19'd18302: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=52;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=842;
 end   
19'd18303: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=41;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=676;
 end   
19'd18304: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=54;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=894;
 end   
19'd18305: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=13;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=248;
 end   
19'd18306: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=62;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=1042;
 end   
19'd18307: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=96;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=1596;
 end   
19'd18308: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=60;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=1030;
 end   
19'd18309: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=4;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=572;
 end   
19'd18310: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=99;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=2327;
 end   
19'd18311: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=36;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=1216;
 end   
19'd18312: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=80;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=2094;
 end   
19'd18313: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=98;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=1718;
 end   
19'd18314: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=32;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=1522;
 end   
19'd18315: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=87;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=2901;
 end   
19'd18316: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=84;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=2290;
 end   
19'd18317: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd18459: begin  
rid<=1;
end
19'd18460: begin  
end
19'd18461: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd18462: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd18463: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd18464: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd18465: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd18466: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd18467: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd18468: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd18469: begin  
rid<=0;
end
19'd18601: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=82;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4865;
 end   
19'd18602: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=49;
   mapp<=70;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4292;
 end   
19'd18603: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=23;
   mapp<=41;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4423;
 end   
19'd18604: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=58;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1589;
 end   
19'd18605: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=5;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5435;
 end   
19'd18606: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=21;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=10762;
 end   
19'd18607: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=95;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=8006;
 end   
19'd18608: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=96;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd18609: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd18610: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=58;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=19345;
 end   
19'd18611: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=77;
   mapp<=78;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=14751;
 end   
19'd18612: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=50;
   mapp<=79;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=11160;
 end   
19'd18613: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=7;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=10796;
 end   
19'd18614: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=29;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=21520;
 end   
19'd18615: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=81;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=30652;
 end   
19'd18616: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=95;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=27504;
 end   
19'd18617: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=78;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd18618: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=76;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd18619: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd18761: begin  
rid<=1;
end
19'd18762: begin  
end
19'd18763: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd18764: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd18765: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd18766: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd18767: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd18768: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd18769: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd18770: begin  
rid<=0;
end
19'd18901: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=65;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5460;
 end   
19'd18902: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=93;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7822;
 end   
19'd18903: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=8;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=692;
 end   
19'd18904: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=72;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6078;
 end   
19'd18905: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=43;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3652;
 end   
19'd18906: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=29;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=2486;
 end   
19'd18907: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=14;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=1236;
 end   
19'd18908: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=68;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=5782;
 end   
19'd18909: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=55;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=4700;
 end   
19'd18910: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=91;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=7734;
 end   
19'd18911: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=73;
   mapp<=0;
   pp<=100;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[10]<=6232;
 end   
19'd18912: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=48;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=6516;
 end   
19'd18913: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=51;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8944;
 end   
19'd18914: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=86;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=2584;
 end   
19'd18915: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=44;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=7046;
 end   
19'd18916: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=46;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=4664;
 end   
19'd18917: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=77;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=4180;
 end   
19'd18918: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=17;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=1610;
 end   
19'd18919: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=29;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=6420;
 end   
19'd18920: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=16;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=5052;
 end   
19'd18921: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=74;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=9362;
 end   
19'd18922: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=91;
   mapp<=0;
   pp<=100;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[10]<=8234;
 end   
19'd18923: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd19065: begin  
rid<=1;
end
19'd19066: begin  
end
19'd19067: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd19068: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd19069: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd19070: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd19071: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd19072: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd19073: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd19074: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd19075: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd19076: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd19077: begin  
check0<=expctdoutput[10]-outcheck0;
end
19'd19078: begin  
rid<=0;
end
19'd19201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=49;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11975;
 end   
19'd19202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=57;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11624;
 end   
19'd19203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=40;
   mapp<=91;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10737;
 end   
19'd19204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=52;
   mapp<=15;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=11716;
 end   
19'd19205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=36;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=14746;
 end   
19'd19206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=51;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=13783;
 end   
19'd19207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=87;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=12947;
 end   
19'd19208: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=26;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=13282;
 end   
19'd19209: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd19210: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=55;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd19211: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=83;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd19212: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=65;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=30112;
 end   
19'd19213: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=13;
   mapp<=80;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=30362;
 end   
19'd19214: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=61;
   mapp<=97;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=35347;
 end   
19'd19215: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=78;
   mapp<=65;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=35454;
 end   
19'd19216: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=78;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=32913;
 end   
19'd19217: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=78;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=28437;
 end   
19'd19218: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=40;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=25071;
 end   
19'd19219: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=11;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=26991;
 end   
19'd19220: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=47;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd19221: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=45;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd19222: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd19223: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd19365: begin  
rid<=1;
end
19'd19366: begin  
end
19'd19367: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd19368: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd19369: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd19370: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd19371: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd19372: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd19373: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd19374: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd19375: begin  
rid<=0;
end
19'd19501: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=49;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2450;
 end   
19'd19502: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=33;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1660;
 end   
19'd19503: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=65;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3270;
 end   
19'd19504: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=14;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=730;
 end   
19'd19505: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=7;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=3024;
 end   
19'd19506: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=32;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=4284;
 end   
19'd19507: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=96;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=11142;
 end   
19'd19508: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=67;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6224;
 end   
19'd19509: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd19651: begin  
rid<=1;
end
19'd19652: begin  
end
19'd19653: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd19654: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd19655: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd19656: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd19657: begin  
rid<=0;
end
19'd19801: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=46;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=24454;
 end   
19'd19802: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=76;
   mapp<=41;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=20455;
 end   
19'd19803: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=59;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd19804: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=89;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd19805: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=22;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd19806: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=66;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd19807: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=86;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd19808: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=55;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd19809: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=28;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd19810: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=14;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd19811: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd19812: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=52;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=51195;
 end   
19'd19813: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=21;
   mapp<=53;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=39795;
 end   
19'd19814: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=96;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd19815: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=81;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd19816: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=21;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd19817: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=55;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd19818: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=47;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd19819: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=24;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd19820: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=18;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd19821: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=35;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd19822: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd19823: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd19965: begin  
rid<=1;
end
19'd19966: begin  
end
19'd19967: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd19968: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd19969: begin  
rid<=0;
end
19'd20101: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=53;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7873;
 end   
19'd20102: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=22;
   mapp<=98;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7920;
 end   
19'd20103: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=35;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd20104: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=43;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd20105: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=47;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17081;
 end   
19'd20106: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=80;
   mapp<=53;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18834;
 end   
19'd20107: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=26;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd20108: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=78;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd20109: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd20251: begin  
rid<=1;
end
19'd20252: begin  
end
19'd20253: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd20254: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd20255: begin  
rid<=0;
end
19'd20401: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=73;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=18750;
 end   
19'd20402: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=61;
   mapp<=99;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=17663;
 end   
19'd20403: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=45;
   mapp<=55;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=18060;
 end   
19'd20404: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=73;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd20405: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=74;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd20406: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=50;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd20407: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=53;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd20408: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=65;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=34476;
 end   
19'd20409: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=72;
   mapp<=87;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=37425;
 end   
19'd20410: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=29;
   mapp<=99;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=32887;
 end   
19'd20411: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=81;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd20412: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=12;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd20413: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=76;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd20414: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=81;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd20415: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd20557: begin  
rid<=1;
end
19'd20558: begin  
end
19'd20559: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd20560: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd20561: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd20562: begin  
rid<=0;
end
19'd20701: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=93;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=20029;
 end   
19'd20702: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=6;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=14456;
 end   
19'd20703: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=78;
   mapp<=72;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=21229;
 end   
19'd20704: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=48;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd20705: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=6;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd20706: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=71;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd20707: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=66;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd20708: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd20709: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd20710: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=78;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=40384;
 end   
19'd20711: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=17;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=33034;
 end   
19'd20712: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=15;
   mapp<=20;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=33992;
 end   
19'd20713: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=26;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd20714: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=84;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd20715: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=68;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd20716: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=6;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd20717: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd20718: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd20719: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd20861: begin  
rid<=1;
end
19'd20862: begin  
end
19'd20863: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd20864: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd20865: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd20866: begin  
rid<=0;
end
19'd21001: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=99;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9432;
 end   
19'd21002: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=85;
   mapp<=90;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9280;
 end   
19'd21003: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=86;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10478;
 end   
19'd21004: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=99;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3612;
 end   
19'd21005: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=20;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1300;
 end   
19'd21006: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=10;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6620;
 end   
19'd21007: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=71;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=2508;
 end   
19'd21008: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=13;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=1654;
 end   
19'd21009: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=15;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd21010: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=80;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16790;
 end   
19'd21011: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=31;
   mapp<=18;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=13121;
 end   
19'd21012: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=67;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=17739;
 end   
19'd21013: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=87;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=11799;
 end   
19'd21014: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=44;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=6588;
 end   
19'd21015: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=86;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=14056;
 end   
19'd21016: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=7;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=4183;
 end   
19'd21017: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=60;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=7240;
 end   
19'd21018: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=27;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd21019: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd21161: begin  
rid<=1;
end
19'd21162: begin  
end
19'd21163: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd21164: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd21165: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd21166: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd21167: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd21168: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd21169: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd21170: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd21171: begin  
rid<=0;
end
19'd21301: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=93;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13387;
 end   
19'd21302: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=85;
   mapp<=71;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7805;
 end   
19'd21303: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=37;
   mapp<=68;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2997;
 end   
19'd21304: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=11;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6122;
 end   
19'd21305: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=4;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6123;
 end   
19'd21306: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=77;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=9104;
 end   
19'd21307: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=6;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=6696;
 end   
19'd21308: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=68;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=6052;
 end   
19'd21309: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=22;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd21310: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=13;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd21311: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=19118;
 end   
19'd21312: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=88;
   mapp<=42;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=13408;
 end   
19'd21313: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=55;
   mapp<=37;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=8474;
 end   
19'd21314: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=89;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=11093;
 end   
19'd21315: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=47;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=12966;
 end   
19'd21316: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=81;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=16118;
 end   
19'd21317: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=93;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=13443;
 end   
19'd21318: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=84;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=11963;
 end   
19'd21319: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=87;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd21320: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=61;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd21321: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd21463: begin  
rid<=1;
end
19'd21464: begin  
end
19'd21465: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd21466: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd21467: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd21468: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd21469: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd21470: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd21471: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd21472: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd21473: begin  
rid<=0;
end
19'd21601: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=82;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=82;
 end   
19'd21602: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=65;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=3137;
 end   
19'd21603: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd21745: begin  
rid<=1;
end
19'd21746: begin  
end
19'd21747: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd21748: begin  
rid<=0;
end
19'd21901: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=6;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=20452;
 end   
19'd21902: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=56;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=21075;
 end   
19'd21903: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=43;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd21904: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=93;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd21905: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=80;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd21906: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=80;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd21907: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd21908: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=68;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=33200;
 end   
19'd21909: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=40;
   mapp<=11;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=32375;
 end   
19'd21910: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=31;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd21911: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=33;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd21912: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=79;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd21913: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=63;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd21914: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd21915: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd22057: begin  
rid<=1;
end
19'd22058: begin  
end
19'd22059: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd22060: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd22061: begin  
rid<=0;
end
19'd22201: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=80;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2880;
 end   
19'd22202: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7610;
 end   
19'd22203: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=65;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5220;
 end   
19'd22204: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=74;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5950;
 end   
19'd22205: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=20;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1640;
 end   
19'd22206: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=35;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=2850;
 end   
19'd22207: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=56;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7136;
 end   
19'd22208: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=55;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=10690;
 end   
19'd22209: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=25;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=6620;
 end   
19'd22210: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=71;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=9926;
 end   
19'd22211: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=8;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=2088;
 end   
19'd22212: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=59;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=6154;
 end   
19'd22213: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd22355: begin  
rid<=1;
end
19'd22356: begin  
end
19'd22357: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd22358: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd22359: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd22360: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd22361: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd22362: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd22363: begin  
rid<=0;
end
19'd22501: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=85;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2905;
 end   
19'd22502: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=62;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8060;
 end   
19'd22503: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=75;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10239;
 end   
19'd22504: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd22505: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=8;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=6425;
 end   
19'd22506: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=80;
   mapp<=36;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=16108;
 end   
19'd22507: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=97;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=11175;
 end   
19'd22508: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd22509: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd22651: begin  
rid<=1;
end
19'd22652: begin  
end
19'd22653: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd22654: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd22655: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd22656: begin  
rid<=0;
end
19'd22801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=97;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=18289;
 end   
19'd22802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=80;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15318;
 end   
19'd22803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=35;
   mapp<=40;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=17956;
 end   
19'd22804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=72;
   mapp<=46;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=14893;
 end   
19'd22805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=74;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=15385;
 end   
19'd22806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=7;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd22807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=55;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd22808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=66;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd22809: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=41;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd22810: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd22811: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=12;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=29939;
 end   
19'd22812: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=36;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=28271;
 end   
19'd22813: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=55;
   mapp<=15;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=32027;
 end   
19'd22814: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=62;
   mapp<=96;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=26143;
 end   
19'd22815: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=43;
   mapp<=25;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=24883;
 end   
19'd22816: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=42;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd22817: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=21;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd22818: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=22;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd22819: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd22820: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=48;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd22821: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd22963: begin  
rid<=1;
end
19'd22964: begin  
end
19'd22965: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd22966: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd22967: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd22968: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd22969: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd22970: begin  
rid<=0;
end
19'd23101: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=35;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=595;
 end   
19'd23102: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=14;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=500;
 end   
19'd23103: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=50;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1770;
 end   
19'd23104: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=90;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3180;
 end   
19'd23105: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=40;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=2955;
 end   
19'd23106: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=69;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=3260;
 end   
19'd23107: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=95;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=5570;
 end   
19'd23108: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=3;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=3300;
 end   
19'd23109: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd23251: begin  
rid<=1;
end
19'd23252: begin  
end
19'd23253: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd23254: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd23255: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd23256: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd23257: begin  
rid<=0;
end
19'd23401: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=61;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7676;
 end   
19'd23402: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=81;
   mapp<=91;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5147;
 end   
19'd23403: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=52;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5103;
 end   
19'd23404: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=53;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3298;
 end   
19'd23405: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=33;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2844;
 end   
19'd23406: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=29;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=8112;
 end   
19'd23407: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=87;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=4317;
 end   
19'd23408: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=42;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=5103;
 end   
19'd23409: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=53;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=7898;
 end   
19'd23410: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=83;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=2325;
 end   
19'd23411: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=20;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd23412: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=44;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=9426;
 end   
19'd23413: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=63;
   mapp<=18;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=6551;
 end   
19'd23414: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=29;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=6445;
 end   
19'd23415: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=52;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=5178;
 end   
19'd23416: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=64;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=4982;
 end   
19'd23417: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=69;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=10338;
 end   
19'd23418: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=70;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=5387;
 end   
19'd23419: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=5;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=6019;
 end   
19'd23420: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=47;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=10248;
 end   
19'd23421: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=94;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=5207;
 end   
19'd23422: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=87;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd23423: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd23565: begin  
rid<=1;
end
19'd23566: begin  
end
19'd23567: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd23568: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd23569: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd23570: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd23571: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd23572: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd23573: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd23574: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd23575: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd23576: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd23577: begin  
rid<=0;
end
19'd23701: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=71;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=19586;
 end   
19'd23702: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=45;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=23267;
 end   
19'd23703: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=21;
   mapp<=79;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=23490;
 end   
19'd23704: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=70;
   mapp<=90;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=24595;
 end   
19'd23705: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=83;
   mapp<=88;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=23886;
 end   
19'd23706: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=89;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd23707: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=55;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd23708: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=78;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd23709: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=79;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd23710: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=6;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd23711: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=35;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=49018;
 end   
19'd23712: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=79;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=47435;
 end   
19'd23713: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=93;
   mapp<=87;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=44513;
 end   
19'd23714: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=90;
   mapp<=96;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=38877;
 end   
19'd23715: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=62;
   mapp<=33;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=36699;
 end   
19'd23716: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=65;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd23717: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=1;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd23718: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=5;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd23719: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=7;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd23720: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=67;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd23721: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd23863: begin  
rid<=1;
end
19'd23864: begin  
end
19'd23865: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd23866: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd23867: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd23868: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd23869: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd23870: begin  
rid<=0;
end
19'd24001: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=72;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=18434;
 end   
19'd24002: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=63;
   mapp<=57;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=16443;
 end   
19'd24003: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=28;
   mapp<=98;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=16817;
 end   
19'd24004: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=64;
   mapp<=45;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=16635;
 end   
19'd24005: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=1;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd24006: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=23;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd24007: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=90;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd24008: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=4;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd24009: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=1;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd24010: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=27;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd24011: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=97;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd24012: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=45;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=34578;
 end   
19'd24013: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=10;
   mapp<=71;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=30670;
 end   
19'd24014: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=95;
   mapp<=63;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=38922;
 end   
19'd24015: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=41;
   mapp<=1;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=31719;
 end   
19'd24016: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=22;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd24017: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=12;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd24018: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=51;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd24019: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=15;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd24020: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=55;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd24021: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=93;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd24022: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd24023: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd24165: begin  
rid<=1;
end
19'd24166: begin  
end
19'd24167: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd24168: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd24169: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd24170: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd24171: begin  
rid<=0;
end
19'd24301: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=54;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=432;
 end   
19'd24302: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=22;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=186;
 end   
19'd24303: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=7;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=76;
 end   
19'd24304: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=45;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=390;
 end   
19'd24305: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=38;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=344;
 end   
19'd24306: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=44;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=402;
 end   
19'd24307: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=39;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=3942;
 end   
19'd24308: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=54;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=5046;
 end   
19'd24309: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=4;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=436;
 end   
19'd24310: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=23;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=2460;
 end   
19'd24311: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=25;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=2594;
 end   
19'd24312: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=78;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=7422;
 end   
19'd24313: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd24455: begin  
rid<=1;
end
19'd24456: begin  
end
19'd24457: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd24458: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd24459: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd24460: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd24461: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd24462: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd24463: begin  
rid<=0;
end
19'd24601: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=89;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11573;
 end   
19'd24602: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=38;
   mapp<=33;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15255;
 end   
19'd24603: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=63;
   mapp<=23;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=17578;
 end   
19'd24604: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=35;
   mapp<=94;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=19844;
 end   
19'd24605: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=97;
   mapp<=30;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=11999;
 end   
19'd24606: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=46;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=12012;
 end   
19'd24607: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=87;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=15238;
 end   
19'd24608: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd24609: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd24610: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd24611: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd24612: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=61;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17393;
 end   
19'd24613: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=56;
   mapp<=30;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=27135;
 end   
19'd24614: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=6;
   mapp<=24;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=27428;
 end   
19'd24615: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=84;
   mapp<=8;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=29928;
 end   
19'd24616: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=75;
   mapp<=37;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=31543;
 end   
19'd24617: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=74;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=30015;
 end   
19'd24618: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=20;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=28218;
 end   
19'd24619: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd24620: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd24621: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd24622: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd24623: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd24765: begin  
rid<=1;
end
19'd24766: begin  
end
19'd24767: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd24768: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd24769: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd24770: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd24771: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd24772: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd24773: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd24774: begin  
rid<=0;
end
19'd24901: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=79;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12739;
 end   
19'd24902: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=79;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11533;
 end   
19'd24903: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=83;
   mapp<=84;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8591;
 end   
19'd24904: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=67;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6029;
 end   
19'd24905: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=36;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3828;
 end   
19'd24906: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=25;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd24907: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=18;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd24908: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=77;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=18353;
 end   
19'd24909: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=37;
   mapp<=28;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=16514;
 end   
19'd24910: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=91;
   mapp<=19;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15331;
 end   
19'd24911: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=56;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=11901;
 end   
19'd24912: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=95;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=9042;
 end   
19'd24913: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=60;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd24914: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=1;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd24915: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd25057: begin  
rid<=1;
end
19'd25058: begin  
end
19'd25059: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd25060: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd25061: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd25062: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd25063: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd25064: begin  
rid<=0;
end
19'd25201: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=74;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2664;
 end   
19'd25202: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=80;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5930;
 end   
19'd25203: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=75;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5570;
 end   
19'd25204: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=7;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=548;
 end   
19'd25205: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=84;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6256;
 end   
19'd25206: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=29;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=3215;
 end   
19'd25207: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=90;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8540;
 end   
19'd25208: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=76;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=7774;
 end   
19'd25209: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=41;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=1737;
 end   
19'd25210: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=51;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=7735;
 end   
19'd25211: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd25353: begin  
rid<=1;
end
19'd25354: begin  
end
19'd25355: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd25356: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd25357: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd25358: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd25359: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd25360: begin  
rid<=0;
end
19'd25501: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=5;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=37848;
 end   
19'd25502: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=76;
   mapp<=91;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=35691;
 end   
19'd25503: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=79;
   mapp<=89;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=31297;
 end   
19'd25504: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=95;
   mapp<=87;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=33510;
 end   
19'd25505: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=39;
   mapp<=90;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=24095;
 end   
19'd25506: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=68;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd25507: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=98;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd25508: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd25509: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd25510: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd25511: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd25512: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=78;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=54477;
 end   
19'd25513: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=91;
   mapp<=39;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=48272;
 end   
19'd25514: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=23;
   mapp<=15;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=41389;
 end   
19'd25515: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=43;
   mapp<=21;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=51620;
 end   
19'd25516: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=34;
   mapp<=93;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=45141;
 end   
19'd25517: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=43;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd25518: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=49;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd25519: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd25520: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd25521: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd25522: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd25523: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd25665: begin  
rid<=1;
end
19'd25666: begin  
end
19'd25667: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd25668: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd25669: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd25670: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd25671: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd25672: begin  
rid<=0;
end
19'd25801: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=16;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14463;
 end   
19'd25802: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=90;
   mapp<=41;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15625;
 end   
19'd25803: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=62;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd25804: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=35;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd25805: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=26;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd25806: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=10;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd25807: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=77;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd25808: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd25809: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=66;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=32420;
 end   
19'd25810: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=60;
   mapp<=60;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=39675;
 end   
19'd25811: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=38;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd25812: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=88;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd25813: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=11;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd25814: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=45;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd25815: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=67;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd25816: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd25817: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd25959: begin  
rid<=1;
end
19'd25960: begin  
end
19'd25961: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd25962: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd25963: begin  
rid<=0;
end
19'd26101: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=3;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9844;
 end   
19'd26102: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=48;
   mapp<=42;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12051;
 end   
19'd26103: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=51;
   mapp<=63;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8655;
 end   
19'd26104: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=70;
   mapp<=47;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=10400;
 end   
19'd26105: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=36;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd26106: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=58;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd26107: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd26108: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd26109: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd26110: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=95;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=24962;
 end   
19'd26111: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=44;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=23395;
 end   
19'd26112: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=91;
   mapp<=5;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=23633;
 end   
19'd26113: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=3;
   mapp<=31;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=23420;
 end   
19'd26114: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=88;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd26115: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=15;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd26116: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd26117: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd26118: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd26119: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd26261: begin  
rid<=1;
end
19'd26262: begin  
end
19'd26263: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd26264: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd26265: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd26266: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd26267: begin  
rid<=0;
end
19'd26401: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=75;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14949;
 end   
19'd26402: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=42;
   mapp<=91;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11095;
 end   
19'd26403: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=69;
   mapp<=83;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12044;
 end   
19'd26404: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=33;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=14223;
 end   
19'd26405: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=54;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=19962;
 end   
19'd26406: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=78;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=19221;
 end   
19'd26407: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=85;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=17175;
 end   
19'd26408: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=57;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=17866;
 end   
19'd26409: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=33;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd26410: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=93;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd26411: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=90;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd26412: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=71;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=19518;
 end   
19'd26413: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=11;
   mapp<=50;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=17784;
 end   
19'd26414: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=90;
   mapp<=33;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=16843;
 end   
19'd26415: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=38;
   mapp<=22;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=19335;
 end   
19'd26416: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=41;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=25680;
 end   
19'd26417: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=58;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=24737;
 end   
19'd26418: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=47;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=23568;
 end   
19'd26419: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=52;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=23573;
 end   
19'd26420: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=58;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd26421: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=79;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd26422: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=2;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd26423: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd26565: begin  
rid<=1;
end
19'd26566: begin  
end
19'd26567: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd26568: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd26569: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd26570: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd26571: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd26572: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd26573: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd26574: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd26575: begin  
rid<=0;
end
19'd26701: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=95;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2746;
 end   
19'd26702: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=35;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1966;
 end   
19'd26703: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=8;
   mapp<=22;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5108;
 end   
19'd26704: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=61;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd26705: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=42;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd26706: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=78;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=19252;
 end   
19'd26707: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=42;
   mapp<=99;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=15165;
 end   
19'd26708: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=57;
   mapp<=88;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=18661;
 end   
19'd26709: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=41;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd26710: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=47;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd26711: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd26853: begin  
rid<=1;
end
19'd26854: begin  
end
19'd26855: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd26856: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd26857: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd26858: begin  
rid<=0;
end
19'd27001: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=13;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1040;
 end   
19'd27002: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=64;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5130;
 end   
19'd27003: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=10;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=820;
 end   
19'd27004: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=61;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4910;
 end   
19'd27005: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=85;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6840;
 end   
19'd27006: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=73;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=5890;
 end   
19'd27007: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=4;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=380;
 end   
19'd27008: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=62;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=5030;
 end   
19'd27009: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=3;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=320;
 end   
19'd27010: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=2;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=250;
 end   
19'd27011: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=69;
   mapp<=0;
   pp<=100;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[10]<=5620;
 end   
19'd27012: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=29;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=2606;
 end   
19'd27013: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=52;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=7938;
 end   
19'd27014: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=74;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=4816;
 end   
19'd27015: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=49;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=7556;
 end   
19'd27016: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=30;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=8460;
 end   
19'd27017: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=44;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=8266;
 end   
19'd27018: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=44;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=2756;
 end   
19'd27019: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=49;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=7676;
 end   
19'd27020: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=18;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=1292;
 end   
19'd27021: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=65;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=3760;
 end   
19'd27022: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=63;
   mapp<=0;
   pp<=100;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[10]<=9022;
 end   
19'd27023: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd27165: begin  
rid<=1;
end
19'd27166: begin  
end
19'd27167: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd27168: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd27169: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd27170: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd27171: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd27172: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd27173: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd27174: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd27175: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd27176: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd27177: begin  
check0<=expctdoutput[10]-outcheck0;
end
19'd27178: begin  
rid<=0;
end
19'd27301: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=98;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=18137;
 end   
19'd27302: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=3;
   mapp<=31;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11251;
 end   
19'd27303: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=52;
   mapp<=47;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=19215;
 end   
19'd27304: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=79;
   mapp<=11;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=21712;
 end   
19'd27305: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=53;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd27306: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=43;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd27307: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=22;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd27308: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd27309: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=63;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd27310: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=51;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=34217;
 end   
19'd27311: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=80;
   mapp<=50;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=23911;
 end   
19'd27312: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=77;
   mapp<=22;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=29025;
 end   
19'd27313: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=16;
   mapp<=40;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=33153;
 end   
19'd27314: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=76;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd27315: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=78;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd27316: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=20;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd27317: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=15;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd27318: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=48;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd27319: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd27461: begin  
rid<=1;
end
19'd27462: begin  
end
19'd27463: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd27464: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd27465: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd27466: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd27467: begin  
rid<=0;
end
19'd27601: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=62;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7430;
 end   
19'd27602: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=2;
   mapp<=57;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5274;
 end   
19'd27603: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=62;
   mapp<=83;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9140;
 end   
19'd27604: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=20;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd27605: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd27606: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=86;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16443;
 end   
19'd27607: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=88;
   mapp<=73;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=9148;
 end   
19'd27608: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=17;
   mapp<=41;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=14527;
 end   
19'd27609: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=17;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd27610: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=92;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd27611: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd27753: begin  
rid<=1;
end
19'd27754: begin  
end
19'd27755: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd27756: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd27757: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd27758: begin  
rid<=0;
end
19'd27901: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=19;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7423;
 end   
19'd27902: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=81;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd27903: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=3;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd27904: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=30;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd27905: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=30;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16555;
 end   
19'd27906: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=72;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd27907: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=64;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd27908: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=7;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd27909: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd28051: begin  
rid<=1;
end
19'd28052: begin  
end
19'd28053: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd28054: begin  
rid<=0;
end
19'd28201: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=33;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=22812;
 end   
19'd28202: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=37;
   mapp<=90;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=24438;
 end   
19'd28203: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=93;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd28204: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=30;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd28205: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=74;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd28206: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=93;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd28207: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=82;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd28208: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=3;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd28209: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd28210: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=40;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=47896;
 end   
19'd28211: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=3;
   mapp<=90;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=46717;
 end   
19'd28212: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=66;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd28213: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=83;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd28214: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=61;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd28215: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=59;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd28216: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=45;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd28217: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=86;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd28218: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd28219: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd28361: begin  
rid<=1;
end
19'd28362: begin  
end
19'd28363: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd28364: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd28365: begin  
rid<=0;
end
19'd28501: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=83;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4642;
 end   
19'd28502: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=50;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9844;
 end   
19'd28503: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=58;
   mapp<=9;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9450;
 end   
19'd28504: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=21;
   mapp<=97;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=12219;
 end   
19'd28505: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=75;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=11025;
 end   
19'd28506: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=81;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd28507: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=87;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd28508: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=71;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd28509: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=38;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12887;
 end   
19'd28510: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=99;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=14480;
 end   
19'd28511: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=30;
   mapp<=4;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=18566;
 end   
19'd28512: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=61;
   mapp<=79;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=22488;
 end   
19'd28513: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=18;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=15458;
 end   
19'd28514: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=5;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd28515: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=40;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd28516: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=28;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd28517: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd28659: begin  
rid<=1;
end
19'd28660: begin  
end
19'd28661: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd28662: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd28663: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd28664: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd28665: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd28666: begin  
rid<=0;
end
19'd28801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=93;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=29066;
 end   
19'd28802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=96;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd28803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=61;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd28804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=46;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd28805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=38;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd28806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=70;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd28807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=38;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd28808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=33;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=42800;
 end   
19'd28809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=55;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd28810: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=65;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd28811: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=26;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd28812: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=1;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd28813: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=34;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd28814: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=59;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd28815: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd28957: begin  
rid<=1;
end
19'd28958: begin  
end
19'd28959: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd28960: begin  
rid<=0;
end
19'd29101: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=27;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10987;
 end   
19'd29102: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=98;
   mapp<=92;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11608;
 end   
19'd29103: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=93;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5765;
 end   
19'd29104: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=33;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4547;
 end   
19'd29105: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=37;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1333;
 end   
19'd29106: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=3;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=8951;
 end   
19'd29107: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=90;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=3568;
 end   
19'd29108: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=11;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=9579;
 end   
19'd29109: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=94;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=9282;
 end   
19'd29110: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd29111: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=36;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=18943;
 end   
19'd29112: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=99;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=21157;
 end   
19'd29113: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=79;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=13262;
 end   
19'd29114: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=47;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=11090;
 end   
19'd29115: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=49;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=6166;
 end   
19'd29116: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=31;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=16898;
 end   
19'd29117: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=69;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=13477;
 end   
19'd29118: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=75;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=21981;
 end   
19'd29119: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=98;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=17661;
 end   
19'd29120: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd29121: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd29263: begin  
rid<=1;
end
19'd29264: begin  
end
19'd29265: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd29266: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd29267: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd29268: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd29269: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd29270: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd29271: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd29272: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd29273: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd29274: begin  
rid<=0;
end
19'd29401: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=67;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8614;
 end   
19'd29402: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=16;
   mapp<=54;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7766;
 end   
19'd29403: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=93;
   mapp<=61;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12556;
 end   
19'd29404: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd29405: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd29406: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=84;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=18573;
 end   
19'd29407: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=92;
   mapp<=66;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18722;
 end   
19'd29408: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=67;
   mapp<=53;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=19285;
 end   
19'd29409: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd29410: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd29411: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd29553: begin  
rid<=1;
end
19'd29554: begin  
end
19'd29555: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd29556: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd29557: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd29558: begin  
rid<=0;
end
19'd29701: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=4;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13451;
 end   
19'd29702: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=99;
   mapp<=11;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11057;
 end   
19'd29703: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=74;
   mapp<=14;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=13486;
 end   
19'd29704: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=95;
   mapp<=90;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=13721;
 end   
19'd29705: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=6;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd29706: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=58;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd29707: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd29708: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=58;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd29709: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=9;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd29710: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=26;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=25024;
 end   
19'd29711: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=89;
   mapp<=47;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=29785;
 end   
19'd29712: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=3;
   mapp<=40;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=28235;
 end   
19'd29713: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=66;
   mapp<=18;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=35008;
 end   
19'd29714: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=12;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd29715: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=40;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd29716: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd29717: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=76;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd29718: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=95;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd29719: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd29861: begin  
rid<=1;
end
19'd29862: begin  
end
19'd29863: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd29864: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd29865: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd29866: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd29867: begin  
rid<=0;
end
19'd30001: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=81;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4131;
 end   
19'd30002: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=9;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=739;
 end   
19'd30003: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=87;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7067;
 end   
19'd30004: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=83;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6753;
 end   
19'd30005: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=85;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6925;
 end   
19'd30006: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=90;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7340;
 end   
19'd30007: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=50;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=4110;
 end   
19'd30008: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=86;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=7036;
 end   
19'd30009: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=55;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=4535;
 end   
19'd30010: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=28;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=4915;
 end   
19'd30011: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=795;
 end   
19'd30012: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=77;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=9223;
 end   
19'd30013: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=62;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=8489;
 end   
19'd30014: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=24;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=7597;
 end   
19'd30015: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=65;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=9160;
 end   
19'd30016: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=72;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=6126;
 end   
19'd30017: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=32;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=7932;
 end   
19'd30018: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=85;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=6915;
 end   
19'd30019: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd30161: begin  
rid<=1;
end
19'd30162: begin  
end
19'd30163: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd30164: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd30165: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd30166: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd30167: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd30168: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd30169: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd30170: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd30171: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd30172: begin  
rid<=0;
end
19'd30301: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=65;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5070;
 end   
19'd30302: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5405;
 end   
19'd30303: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=25;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1645;
 end   
19'd30304: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=21;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=6330;
 end   
19'd30305: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=45;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=6350;
 end   
19'd30306: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=78;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=3283;
 end   
19'd30307: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd30449: begin  
rid<=1;
end
19'd30450: begin  
end
19'd30451: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd30452: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd30453: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd30454: begin  
rid<=0;
end
19'd30601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=1;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2728;
 end   
19'd30602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=37;
   mapp<=73;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1341;
 end   
19'd30603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=34;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1941;
 end   
19'd30604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=51;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=2856;
 end   
19'd30605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=75;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1447;
 end   
19'd30606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=36;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=1344;
 end   
19'd30607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd30608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=45;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=9246;
 end   
19'd30609: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=82;
   mapp<=74;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12051;
 end   
19'd30610: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=90;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=10583;
 end   
19'd30611: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=56;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=11198;
 end   
19'd30612: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=71;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=11202;
 end   
19'd30613: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=80;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=7814;
 end   
19'd30614: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd30615: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd30757: begin  
rid<=1;
end
19'd30758: begin  
end
19'd30759: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd30760: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd30761: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd30762: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd30763: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd30764: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd30765: begin  
rid<=0;
end
19'd30901: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=3;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16469;
 end   
19'd30902: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=31;
   mapp<=12;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=14753;
 end   
19'd30903: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=15;
   mapp<=37;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=15489;
 end   
19'd30904: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=39;
   mapp<=98;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=14978;
 end   
19'd30905: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=58;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd30906: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=29;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd30907: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=45;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd30908: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=94;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd30909: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd30910: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd30911: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd30912: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=8;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=39249;
 end   
19'd30913: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=3;
   mapp<=45;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=34531;
 end   
19'd30914: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=77;
   mapp<=72;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=36344;
 end   
19'd30915: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=25;
   mapp<=75;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=36901;
 end   
19'd30916: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=34;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd30917: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=1;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd30918: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=78;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd30919: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=82;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd30920: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd30921: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd30922: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd30923: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd31065: begin  
rid<=1;
end
19'd31066: begin  
end
19'd31067: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd31068: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd31069: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd31070: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd31071: begin  
rid<=0;
end
19'd31201: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=75;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6786;
 end   
19'd31202: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=24;
   mapp<=39;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3847;
 end   
19'd31203: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=38;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3374;
 end   
19'd31204: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=21;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=2229;
 end   
19'd31205: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=26;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3502;
 end   
19'd31206: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=63;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6623;
 end   
19'd31207: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd31208: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=84;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=13590;
 end   
19'd31209: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=16;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=4823;
 end   
19'd31210: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=61;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=9490;
 end   
19'd31211: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=62;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=7469;
 end   
19'd31212: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=2;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=4438;
 end   
19'd31213: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=48;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=12175;
 end   
19'd31214: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd31215: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd31357: begin  
rid<=1;
end
19'd31358: begin  
end
19'd31359: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd31360: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd31361: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd31362: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd31363: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd31364: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd31365: begin  
rid<=0;
end
19'd31501: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=44;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9048;
 end   
19'd31502: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=59;
   mapp<=84;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7261;
 end   
19'd31503: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=21;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6845;
 end   
19'd31504: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=58;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd31505: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=77;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=13651;
 end   
19'd31506: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=19;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=11954;
 end   
19'd31507: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=57;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=12084;
 end   
19'd31508: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=41;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd31509: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd31651: begin  
rid<=1;
end
19'd31652: begin  
end
19'd31653: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd31654: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd31655: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd31656: begin  
rid<=0;
end
19'd31801: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=41;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3292;
 end   
19'd31802: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=15;
   mapp<=15;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4825;
 end   
19'd31803: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=15;
   mapp<=72;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6720;
 end   
19'd31804: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=36;
   mapp<=29;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5961;
 end   
19'd31805: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=57;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3744;
 end   
19'd31806: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=59;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7848;
 end   
19'd31807: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd31808: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=52;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd31809: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=93;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd31810: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=98;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=11156;
 end   
19'd31811: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=24;
   mapp<=29;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=10948;
 end   
19'd31812: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=24;
   mapp<=48;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=13729;
 end   
19'd31813: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=74;
   mapp<=27;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=15058;
 end   
19'd31814: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=33;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=11276;
 end   
19'd31815: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=85;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=17469;
 end   
19'd31816: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd31817: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd31818: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd31819: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd31961: begin  
rid<=1;
end
19'd31962: begin  
end
19'd31963: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd31964: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd31965: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd31966: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd31967: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd31968: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd31969: begin  
rid<=0;
end
19'd32101: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4011;
 end   
19'd32102: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=24;
   mapp<=78;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8467;
 end   
19'd32103: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=93;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd32104: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd32105: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=7;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=10430;
 end   
19'd32106: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=77;
   mapp<=12;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=19184;
 end   
19'd32107: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=84;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd32108: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd32109: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd32251: begin  
rid<=1;
end
19'd32252: begin  
end
19'd32253: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd32254: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd32255: begin  
rid<=0;
end
19'd32401: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=91;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3094;
 end   
19'd32402: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=21;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=724;
 end   
19'd32403: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=85;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2910;
 end   
19'd32404: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=34;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1186;
 end   
19'd32405: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=90;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3100;
 end   
19'd32406: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=42;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=1478;
 end   
19'd32407: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=98;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=3392;
 end   
19'd32408: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=18;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=4642;
 end   
19'd32409: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=21;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=2530;
 end   
19'd32410: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=24;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=4974;
 end   
19'd32411: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=97;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=9528;
 end   
19'd32412: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=76;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=9636;
 end   
19'd32413: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=54;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=6122;
 end   
19'd32414: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=69;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=9326;
 end   
19'd32415: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd32557: begin  
rid<=1;
end
19'd32558: begin  
end
19'd32559: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd32560: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd32561: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd32562: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd32563: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd32564: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd32565: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd32566: begin  
rid<=0;
end
19'd32701: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=2;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2770;
 end   
19'd32702: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=38;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd32703: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=0;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd32704: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=84;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=10108;
 end   
19'd32705: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=39;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd32706: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=56;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd32707: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd32849: begin  
rid<=1;
end
19'd32850: begin  
end
19'd32851: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd32852: begin  
rid<=0;
end
19'd33001: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=39;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4078;
 end   
19'd33002: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=74;
   mapp<=14;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6994;
 end   
19'd33003: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd33004: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=88;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=6945;
 end   
19'd33005: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=41;
   mapp<=27;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=11584;
 end   
19'd33006: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd33007: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd33149: begin  
rid<=1;
end
19'd33150: begin  
end
19'd33151: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd33152: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd33153: begin  
rid<=0;
end
19'd33301: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=4;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=974;
 end   
19'd33302: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=46;
   mapp<=21;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1278;
 end   
19'd33303: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=56;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd33304: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=8;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=3059;
 end   
19'd33305: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=61;
   mapp<=33;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=2916;
 end   
19'd33306: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=33;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd33307: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd33449: begin  
rid<=1;
end
19'd33450: begin  
end
19'd33451: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd33452: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd33453: begin  
rid<=0;
end
19'd33601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=78;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=21486;
 end   
19'd33602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=87;
   mapp<=42;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=20839;
 end   
19'd33603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=13;
   mapp<=42;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=14291;
 end   
19'd33604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=63;
   mapp<=60;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=16687;
 end   
19'd33605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=91;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd33606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=34;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd33607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=15;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd33608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=56;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd33609: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=61;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd33610: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd33611: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=7;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=37067;
 end   
19'd33612: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=84;
   mapp<=59;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=33879;
 end   
19'd33613: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=51;
   mapp<=51;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=26775;
 end   
19'd33614: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=1;
   mapp<=38;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=33161;
 end   
19'd33615: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=89;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd33616: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=58;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd33617: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=41;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd33618: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=90;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd33619: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=13;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd33620: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd33621: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd33763: begin  
rid<=1;
end
19'd33764: begin  
end
19'd33765: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd33766: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd33767: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd33768: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd33769: begin  
rid<=0;
end
19'd33901: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=66;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=17917;
 end   
19'd33902: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=51;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=20301;
 end   
19'd33903: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=75;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd33904: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=28;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd33905: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=32;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd33906: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=61;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd33907: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=69;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd33908: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=92;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=32319;
 end   
19'd33909: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=70;
   mapp<=29;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=27269;
 end   
19'd33910: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=19;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd33911: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=72;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd33912: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=7;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd33913: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=94;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd33914: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=5;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd33915: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd34057: begin  
rid<=1;
end
19'd34058: begin  
end
19'd34059: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd34060: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd34061: begin  
rid<=0;
end
19'd34201: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=71;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4402;
 end   
19'd34202: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=9;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=649;
 end   
19'd34203: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=7;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=517;
 end   
19'd34204: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=38;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=2728;
 end   
19'd34205: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=60;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4300;
 end   
19'd34206: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=71;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=5091;
 end   
19'd34207: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=66;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7966;
 end   
19'd34208: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=47;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=3751;
 end   
19'd34209: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=14;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=1441;
 end   
19'd34210: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=23;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=4246;
 end   
19'd34211: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=29;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=6214;
 end   
19'd34212: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=89;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=10965;
 end   
19'd34213: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd34355: begin  
rid<=1;
end
19'd34356: begin  
end
19'd34357: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd34358: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd34359: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd34360: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd34361: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd34362: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd34363: begin  
rid<=0;
end
19'd34501: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=39;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5868;
 end   
19'd34502: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=66;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd34503: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=60;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=11587;
 end   
19'd34504: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=53;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd34505: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd34647: begin  
rid<=1;
end
19'd34648: begin  
end
19'd34649: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd34650: begin  
rid<=0;
end
19'd34801: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=66;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=31074;
 end   
19'd34802: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=33;
   mapp<=86;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=29624;
 end   
19'd34803: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=60;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd34804: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=19;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd34805: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=31;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd34806: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=38;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd34807: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=67;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd34808: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=76;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd34809: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=98;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd34810: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=14;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd34811: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd34812: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=93;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=43687;
 end   
19'd34813: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=30;
   mapp<=53;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=43117;
 end   
19'd34814: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=17;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd34815: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=43;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd34816: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=76;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd34817: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=14;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd34818: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=26;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd34819: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=17;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd34820: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=34;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd34821: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=20;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd34822: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd34823: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd34965: begin  
rid<=1;
end
19'd34966: begin  
end
19'd34967: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd34968: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd34969: begin  
rid<=0;
end
19'd35101: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=64;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9262;
 end   
19'd35102: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=75;
   mapp<=54;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5602;
 end   
19'd35103: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=66;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5411;
 end   
19'd35104: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=12;
   mapp<=93;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=11232;
 end   
19'd35105: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=15157;
 end   
19'd35106: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=51;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd35107: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=76;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd35108: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=79;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd35109: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=85;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=24171;
 end   
19'd35110: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=72;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18953;
 end   
19'd35111: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=34;
   mapp<=89;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=19533;
 end   
19'd35112: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=44;
   mapp<=61;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=23672;
 end   
19'd35113: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=61;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=25793;
 end   
19'd35114: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=63;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd35115: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=4;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd35116: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=46;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd35117: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd35259: begin  
rid<=1;
end
19'd35260: begin  
end
19'd35261: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd35262: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd35263: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd35264: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd35265: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd35266: begin  
rid<=0;
end
19'd35401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=18;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3472;
 end   
19'd35402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=11;
   mapp<=30;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6691;
 end   
19'd35403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=92;
   mapp<=23;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7946;
 end   
19'd35404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=64;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6228;
 end   
19'd35405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=74;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5282;
 end   
19'd35406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=46;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=8737;
 end   
19'd35407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd35408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd35409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=69;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12663;
 end   
19'd35410: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=91;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=10992;
 end   
19'd35411: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=23;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15084;
 end   
19'd35412: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=61;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=18718;
 end   
19'd35413: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=91;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=17112;
 end   
19'd35414: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=61;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=15676;
 end   
19'd35415: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd35416: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd35417: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd35559: begin  
rid<=1;
end
19'd35560: begin  
end
19'd35561: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd35562: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd35563: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd35564: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd35565: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd35566: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd35567: begin  
rid<=0;
end
19'd35701: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=14;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=238;
 end   
19'd35702: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=95;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1625;
 end   
19'd35703: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=41;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=717;
 end   
19'd35704: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=36;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=642;
 end   
19'd35705: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=67;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1179;
 end   
19'd35706: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=28;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=526;
 end   
19'd35707: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=9;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=715;
 end   
19'd35708: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=73;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=5494;
 end   
19'd35709: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=81;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=5010;
 end   
19'd35710: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=3;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=801;
 end   
19'd35711: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=69;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=4836;
 end   
19'd35712: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=16;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=1374;
 end   
19'd35713: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd35855: begin  
rid<=1;
end
19'd35856: begin  
end
19'd35857: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd35858: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd35859: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd35860: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd35861: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd35862: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd35863: begin  
rid<=0;
end
19'd36001: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=57;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5007;
 end   
19'd36002: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=81;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2554;
 end   
19'd36003: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd36004: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=87;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=11546;
 end   
19'd36005: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=71;
   mapp<=10;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8110;
 end   
19'd36006: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd36007: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd36149: begin  
rid<=1;
end
19'd36150: begin  
end
19'd36151: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd36152: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd36153: begin  
rid<=0;
end
19'd36301: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=71;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6330;
 end   
19'd36302: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=47;
   mapp<=38;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3588;
 end   
19'd36303: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=15;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4476;
 end   
19'd36304: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=92;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6336;
 end   
19'd36305: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=11;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2910;
 end   
19'd36306: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=57;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd36307: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=71;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=10925;
 end   
19'd36308: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=80;
   mapp<=53;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=6108;
 end   
19'd36309: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=40;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=6266;
 end   
19'd36310: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=30;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=10461;
 end   
19'd36311: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=75;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=4345;
 end   
19'd36312: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=20;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd36313: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd36455: begin  
rid<=1;
end
19'd36456: begin  
end
19'd36457: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd36458: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd36459: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd36460: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd36461: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd36462: begin  
rid<=0;
end
19'd36601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=10;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2528;
 end   
19'd36602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=18;
   mapp<=86;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=942;
 end   
19'd36603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=4;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1662;
 end   
19'd36604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=89;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1478;
 end   
19'd36605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=31;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1142;
 end   
19'd36606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=44;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=2074;
 end   
19'd36607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd36608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8192;
 end   
19'd36609: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=96;
   mapp<=59;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=3534;
 end   
19'd36610: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=27;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=2526;
 end   
19'd36611: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=9;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=3302;
 end   
19'd36612: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=19;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=8726;
 end   
19'd36613: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=79;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=3610;
 end   
19'd36614: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd36615: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd36757: begin  
rid<=1;
end
19'd36758: begin  
end
19'd36759: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd36760: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd36761: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd36762: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd36763: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd36764: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd36765: begin  
rid<=0;
end
19'd36901: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=6;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4737;
 end   
19'd36902: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=49;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6502;
 end   
19'd36903: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=54;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8336;
 end   
19'd36904: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=72;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7770;
 end   
19'd36905: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=60;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=10582;
 end   
19'd36906: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=94;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7892;
 end   
19'd36907: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=54;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=4749;
 end   
19'd36908: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=33;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd36909: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=71;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8815;
 end   
19'd36910: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=28;
   mapp<=29;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=9501;
 end   
19'd36911: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=59;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=12239;
 end   
19'd36912: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=41;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=10265;
 end   
19'd36913: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=21;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=14100;
 end   
19'd36914: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=88;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=13854;
 end   
19'd36915: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=66;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=8742;
 end   
19'd36916: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=33;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd36917: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd37059: begin  
rid<=1;
end
19'd37060: begin  
end
19'd37061: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd37062: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd37063: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd37064: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd37065: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd37066: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd37067: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd37068: begin  
rid<=0;
end
19'd37201: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=38;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=18401;
 end   
19'd37202: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=69;
   mapp<=61;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=16302;
 end   
19'd37203: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=83;
   mapp<=60;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12708;
 end   
19'd37204: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=40;
   mapp<=8;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=18788;
 end   
19'd37205: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=95;
   mapp<=82;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=18557;
 end   
19'd37206: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=62;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=21669;
 end   
19'd37207: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=6;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=24372;
 end   
19'd37208: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd37209: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd37210: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd37211: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd37212: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=93;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=31054;
 end   
19'd37213: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=66;
   mapp<=33;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=26748;
 end   
19'd37214: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=51;
   mapp<=9;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=24516;
 end   
19'd37215: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=40;
   mapp<=57;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=32355;
 end   
19'd37216: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=94;
   mapp<=17;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=31937;
 end   
19'd37217: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=34;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=41176;
 end   
19'd37218: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=53;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=42331;
 end   
19'd37219: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd37220: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd37221: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd37222: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd37223: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd37365: begin  
rid<=1;
end
19'd37366: begin  
end
19'd37367: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd37368: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd37369: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd37370: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd37371: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd37372: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd37373: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd37374: begin  
rid<=0;
end
19'd37501: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=51;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9827;
 end   
19'd37502: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=95;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2799;
 end   
19'd37503: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=17;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9148;
 end   
19'd37504: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=92;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=10058;
 end   
19'd37505: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=92;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd37506: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=13;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=13188;
 end   
19'd37507: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=96;
   mapp<=30;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=6651;
 end   
19'd37508: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=10;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=12188;
 end   
19'd37509: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=89;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=14191;
 end   
19'd37510: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=28;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd37511: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd37653: begin  
rid<=1;
end
19'd37654: begin  
end
19'd37655: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd37656: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd37657: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd37658: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd37659: begin  
rid<=0;
end
19'd37801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=82;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6368;
 end   
19'd37802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=69;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3846;
 end   
19'd37803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=20;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4620;
 end   
19'd37804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=93;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7802;
 end   
19'd37805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=92;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6568;
 end   
19'd37806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=62;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=3338;
 end   
19'd37807: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=14;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=1756;
 end   
19'd37808: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=27;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=1538;
 end   
19'd37809: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=7;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=4148;
 end   
19'd37810: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=94;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=4426;
 end   
19'd37811: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=5;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd37812: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=13;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7560;
 end   
19'd37813: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=93;
   mapp<=11;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=5759;
 end   
19'd37814: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=64;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=5485;
 end   
19'd37815: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=3;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=8886;
 end   
19'd37816: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=95;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=8485;
 end   
19'd37817: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=62;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=5035;
 end   
19'd37818: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=81;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=3315;
 end   
19'd37819: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=46;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=2235;
 end   
19'd37820: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=9;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=4793;
 end   
19'd37821: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=48;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=5798;
 end   
19'd37822: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=68;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd37823: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd37965: begin  
rid<=1;
end
19'd37966: begin  
end
19'd37967: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd37968: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd37969: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd37970: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd37971: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd37972: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd37973: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd37974: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd37975: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd37976: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd37977: begin  
rid<=0;
end
19'd38101: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=62;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8533;
 end   
19'd38102: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=27;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7622;
 end   
19'd38103: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=77;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd38104: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=17;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd38105: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=40;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd38106: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=42;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd38107: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=35;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=19549;
 end   
19'd38108: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=30;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=17186;
 end   
19'd38109: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=31;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd38110: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=95;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd38111: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=37;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd38112: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd38113: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd38255: begin  
rid<=1;
end
19'd38256: begin  
end
19'd38257: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd38258: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd38259: begin  
rid<=0;
end
19'd38401: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=80;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2903;
 end   
19'd38402: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=53;
   mapp<=11;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1473;
 end   
19'd38403: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=11;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3762;
 end   
19'd38404: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd38405: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=43;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=6902;
 end   
19'd38406: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=21;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=2376;
 end   
19'd38407: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=85;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=7417;
 end   
19'd38408: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd38409: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd38551: begin  
rid<=1;
end
19'd38552: begin  
end
19'd38553: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd38554: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd38555: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd38556: begin  
rid<=0;
end
19'd38701: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=86;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=18941;
 end   
19'd38702: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=34;
   mapp<=52;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=16554;
 end   
19'd38703: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=48;
   mapp<=75;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=17927;
 end   
19'd38704: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=39;
   mapp<=31;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=19200;
 end   
19'd38705: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=65;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd38706: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=96;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd38707: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=12;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd38708: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd38709: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=52;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd38710: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=31;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd38711: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=82;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=42614;
 end   
19'd38712: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=1;
   mapp<=64;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=38156;
 end   
19'd38713: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=93;
   mapp<=57;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=43476;
 end   
19'd38714: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=99;
   mapp<=48;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=40837;
 end   
19'd38715: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=32;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd38716: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=44;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd38717: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=31;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd38718: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=75;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd38719: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=4;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd38720: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=50;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd38721: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd38863: begin  
rid<=1;
end
19'd38864: begin  
end
19'd38865: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd38866: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd38867: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd38868: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd38869: begin  
rid<=0;
end
19'd39001: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=1;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=38;
 end   
19'd39002: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=23;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=884;
 end   
19'd39003: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=43;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1654;
 end   
19'd39004: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=41;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1588;
 end   
19'd39005: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=80;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3080;
 end   
19'd39006: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=95;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=3660;
 end   
19'd39007: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=18;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=744;
 end   
19'd39008: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=59;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=2312;
 end   
19'd39009: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=63;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=2474;
 end   
19'd39010: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=29;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=850;
 end   
19'd39011: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=88;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=3348;
 end   
19'd39012: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=54;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=3166;
 end   
19'd39013: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=13;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=1952;
 end   
19'd39014: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=79;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=5292;
 end   
19'd39015: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=69;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=5592;
 end   
19'd39016: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=66;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=2592;
 end   
19'd39017: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=79;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=4524;
 end   
19'd39018: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=77;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=4630;
 end   
19'd39019: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd39161: begin  
rid<=1;
end
19'd39162: begin  
end
19'd39163: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd39164: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd39165: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd39166: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd39167: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd39168: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd39169: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd39170: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd39171: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd39172: begin  
rid<=0;
end
19'd39301: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=95;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11109;
 end   
19'd39302: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=97;
   mapp<=92;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11941;
 end   
19'd39303: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=8;
   mapp<=23;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9757;
 end   
19'd39304: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=8;
   mapp<=72;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=12134;
 end   
19'd39305: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=48;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=7639;
 end   
19'd39306: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd39307: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd39308: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd39309: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=5;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=24293;
 end   
19'd39310: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=65;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18632;
 end   
19'd39311: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=23;
   mapp<=65;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=16083;
 end   
19'd39312: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=69;
   mapp<=81;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=14831;
 end   
19'd39313: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=2;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=12807;
 end   
19'd39314: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd39315: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd39316: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd39317: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd39459: begin  
rid<=1;
end
19'd39460: begin  
end
19'd39461: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd39462: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd39463: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd39464: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd39465: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd39466: begin  
rid<=0;
end
19'd39601: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=84;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=420;
 end   
19'd39602: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=78;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=400;
 end   
19'd39603: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=45;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=245;
 end   
19'd39604: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=33;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=1740;
 end   
19'd39605: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=85;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=3800;
 end   
19'd39606: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=245;
 end   
19'd39607: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd39749: begin  
rid<=1;
end
19'd39750: begin  
end
19'd39751: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd39752: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd39753: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd39754: begin  
rid<=0;
end
19'd39901: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=48;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8469;
 end   
19'd39902: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=81;
   mapp<=85;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5403;
 end   
19'd39903: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=32;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5836;
 end   
19'd39904: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=56;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd39905: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=82;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=9361;
 end   
19'd39906: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=1;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=5845;
 end   
19'd39907: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=6;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=8416;
 end   
19'd39908: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=35;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd39909: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd40051: begin  
rid<=1;
end
19'd40052: begin  
end
19'd40053: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd40054: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd40055: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd40056: begin  
rid<=0;
end
19'd40201: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=42;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=18794;
 end   
19'd40202: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=11;
   mapp<=37;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15860;
 end   
19'd40203: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=79;
   mapp<=43;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=19624;
 end   
19'd40204: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=34;
   mapp<=68;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=16870;
 end   
19'd40205: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=12;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd40206: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=93;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd40207: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=30;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd40208: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=61;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd40209: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd40210: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=58;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd40211: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=26;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd40212: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=93;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=37716;
 end   
19'd40213: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=35;
   mapp<=91;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=33358;
 end   
19'd40214: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=24;
   mapp<=43;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=44496;
 end   
19'd40215: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=94;
   mapp<=88;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=40522;
 end   
19'd40216: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=82;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd40217: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=67;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd40218: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=27;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd40219: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=5;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd40220: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=46;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd40221: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=86;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd40222: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd40223: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd40365: begin  
rid<=1;
end
19'd40366: begin  
end
19'd40367: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd40368: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd40369: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd40370: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd40371: begin  
rid<=0;
end
19'd40501: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=77;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7303;
 end   
19'd40502: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=3;
   mapp<=59;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3254;
 end   
19'd40503: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=42;
   mapp<=78;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4378;
 end   
19'd40504: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=56;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5037;
 end   
19'd40505: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=11;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=10739;
 end   
19'd40506: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=25;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=12143;
 end   
19'd40507: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=43;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=9903;
 end   
19'd40508: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=95;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=7158;
 end   
19'd40509: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd40510: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=15;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd40511: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=4;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd40512: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=98;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=10929;
 end   
19'd40513: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=25;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=5651;
 end   
19'd40514: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=13;
   mapp<=41;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=7142;
 end   
19'd40515: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=23;
   mapp<=35;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=8724;
 end   
19'd40516: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=12;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=17732;
 end   
19'd40517: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=18;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=21428;
 end   
19'd40518: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=57;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=21382;
 end   
19'd40519: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=96;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=17202;
 end   
19'd40520: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=39;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd40521: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=86;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd40522: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=94;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd40523: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd40665: begin  
rid<=1;
end
19'd40666: begin  
end
19'd40667: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd40668: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd40669: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd40670: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd40671: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd40672: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd40673: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd40674: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd40675: begin  
rid<=0;
end
19'd40801: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=58;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12343;
 end   
19'd40802: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=47;
   mapp<=11;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=13029;
 end   
19'd40803: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=70;
   mapp<=80;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9875;
 end   
19'd40804: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=90;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd40805: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=73;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd40806: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=27;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd40807: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=50;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=22455;
 end   
19'd40808: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=41;
   mapp<=54;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=21992;
 end   
19'd40809: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=41;
   mapp<=96;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=16228;
 end   
19'd40810: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=46;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd40811: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=25;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd40812: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=13;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd40813: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd40955: begin  
rid<=1;
end
19'd40956: begin  
end
19'd40957: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd40958: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd40959: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd40960: begin  
rid<=0;
end
19'd41101: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=40;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=17714;
 end   
19'd41102: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=79;
   mapp<=3;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=17170;
 end   
19'd41103: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=41;
   mapp<=94;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=13375;
 end   
19'd41104: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=25;
   mapp<=93;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=10443;
 end   
19'd41105: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=34;
   mapp<=67;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=13512;
 end   
19'd41106: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=60;
   mapp<=87;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=22616;
 end   
19'd41107: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd41108: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=7;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd41109: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=21;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd41110: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=92;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd41111: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=93;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd41112: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=11;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=28178;
 end   
19'd41113: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=25;
   mapp<=17;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=28607;
 end   
19'd41114: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=28;
   mapp<=3;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=27743;
 end   
19'd41115: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=78;
   mapp<=43;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=22889;
 end   
19'd41116: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=48;
   mapp<=93;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=23265;
 end   
19'd41117: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=50;
   mapp<=39;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=31690;
 end   
19'd41118: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=92;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd41119: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=44;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd41120: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=54;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd41121: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd41122: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=53;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd41123: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd41265: begin  
rid<=1;
end
19'd41266: begin  
end
19'd41267: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd41268: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd41269: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd41270: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd41271: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd41272: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd41273: begin  
rid<=0;
end
19'd41401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=4;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5503;
 end   
19'd41402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=38;
   mapp<=26;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8850;
 end   
19'd41403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=71;
   mapp<=61;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5827;
 end   
19'd41404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=86;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=10155;
 end   
19'd41405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=5;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6260;
 end   
19'd41406: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=99;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7768;
 end   
19'd41407: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=56;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=7451;
 end   
19'd41408: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=28;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=6211;
 end   
19'd41409: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=67;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=5647;
 end   
19'd41410: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=51;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd41411: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=19;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd41412: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=46;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17306;
 end   
19'd41413: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=93;
   mapp<=66;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=23412;
 end   
19'd41414: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=87;
   mapp<=17;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15334;
 end   
19'd41415: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=21;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=13997;
 end   
19'd41416: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=12;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=13457;
 end   
19'd41417: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=67;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=21147;
 end   
19'd41418: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=99;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=21013;
 end   
19'd41419: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=44;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=16634;
 end   
19'd41420: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=97;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=15016;
 end   
19'd41421: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=1;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd41422: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=28;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd41423: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd41565: begin  
rid<=1;
end
19'd41566: begin  
end
19'd41567: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd41568: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd41569: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd41570: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd41571: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd41572: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd41573: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd41574: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd41575: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd41576: begin  
rid<=0;
end
19'd41701: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=44;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13753;
 end   
19'd41702: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=18;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=18045;
 end   
19'd41703: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=25;
   mapp<=41;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=19948;
 end   
19'd41704: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=19;
   mapp<=96;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=22770;
 end   
19'd41705: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=84;
   mapp<=62;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=23210;
 end   
19'd41706: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=74;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd41707: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=84;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd41708: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=59;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd41709: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=49;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd41710: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=14;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd41711: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=63;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=26880;
 end   
19'd41712: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=51;
   mapp<=3;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=30017;
 end   
19'd41713: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=19;
   mapp<=32;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=28642;
 end   
19'd41714: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=90;
   mapp<=51;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=38781;
 end   
19'd41715: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=17;
   mapp<=37;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=33062;
 end   
19'd41716: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=83;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd41717: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=18;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd41718: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=84;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd41719: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=52;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd41720: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=86;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd41721: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd41863: begin  
rid<=1;
end
19'd41864: begin  
end
19'd41865: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd41866: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd41867: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd41868: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd41869: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd41870: begin  
rid<=0;
end
19'd42001: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=71;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11552;
 end   
19'd42002: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=69;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=14877;
 end   
19'd42003: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=93;
   mapp<=24;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8927;
 end   
19'd42004: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=68;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=11185;
 end   
19'd42005: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=27;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=13918;
 end   
19'd42006: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=48;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=17501;
 end   
19'd42007: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd42008: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd42009: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=92;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=20368;
 end   
19'd42010: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=98;
   mapp<=14;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=24117;
 end   
19'd42011: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=90;
   mapp<=4;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=21397;
 end   
19'd42012: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=84;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=31677;
 end   
19'd42013: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=43;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=28174;
 end   
19'd42014: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=95;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=35689;
 end   
19'd42015: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd42016: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd42017: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd42159: begin  
rid<=1;
end
19'd42160: begin  
end
19'd42161: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd42162: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd42163: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd42164: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd42165: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd42166: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd42167: begin  
rid<=0;
end
19'd42301: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=74;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11495;
 end   
19'd42302: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=14;
   mapp<=74;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10095;
 end   
19'd42303: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=73;
   mapp<=49;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12797;
 end   
19'd42304: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=69;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=10964;
 end   
19'd42305: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=18;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=8141;
 end   
19'd42306: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=65;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=10399;
 end   
19'd42307: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=33;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd42308: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd42309: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=8;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=19675;
 end   
19'd42310: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=49;
   mapp<=52;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18045;
 end   
19'd42311: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=88;
   mapp<=63;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=18058;
 end   
19'd42312: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=45;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=14331;
 end   
19'd42313: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=31;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=9900;
 end   
19'd42314: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=20;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=15404;
 end   
19'd42315: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=6;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd42316: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=71;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd42317: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd42459: begin  
rid<=1;
end
19'd42460: begin  
end
19'd42461: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd42462: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd42463: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd42464: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd42465: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd42466: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd42467: begin  
rid<=0;
end
19'd42601: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=22;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6743;
 end   
19'd42602: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=23;
   mapp<=57;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11394;
 end   
19'd42603: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=6;
   mapp<=47;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11195;
 end   
19'd42604: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=6;
   mapp<=82;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=13711;
 end   
19'd42605: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=89;
   mapp<=38;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=15565;
 end   
19'd42606: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=56;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd42607: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=45;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd42608: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=51;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd42609: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd42610: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=6;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17728;
 end   
19'd42611: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=10;
   mapp<=50;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=24055;
 end   
19'd42612: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=13;
   mapp<=97;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=27236;
 end   
19'd42613: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=51;
   mapp<=36;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=28176;
 end   
19'd42614: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=80;
   mapp<=91;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=28947;
 end   
19'd42615: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=44;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd42616: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=43;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd42617: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=41;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd42618: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=45;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd42619: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd42761: begin  
rid<=1;
end
19'd42762: begin  
end
19'd42763: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd42764: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd42765: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd42766: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd42767: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd42768: begin  
rid<=0;
end
19'd42901: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=24;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5395;
 end   
19'd42902: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=4;
   mapp<=14;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2988;
 end   
19'd42903: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=56;
   mapp<=85;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4318;
 end   
19'd42904: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=17;
   mapp<=27;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5222;
 end   
19'd42905: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=27;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3437;
 end   
19'd42906: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=55;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=9499;
 end   
19'd42907: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=2;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=9700;
 end   
19'd42908: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=86;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=11915;
 end   
19'd42909: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=68;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd42910: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=98;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd42911: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=79;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd42912: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=75;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16976;
 end   
19'd42913: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=10;
   mapp<=89;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=19748;
 end   
19'd42914: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=32;
   mapp<=58;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=22659;
 end   
19'd42915: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=89;
   mapp<=90;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=18725;
 end   
19'd42916: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=96;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=11619;
 end   
19'd42917: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=50;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=15003;
 end   
19'd42918: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=12;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=19952;
 end   
19'd42919: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=22;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=22154;
 end   
19'd42920: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=29;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd42921: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=72;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd42922: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=36;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd42923: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd43065: begin  
rid<=1;
end
19'd43066: begin  
end
19'd43067: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd43068: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd43069: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd43070: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd43071: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd43072: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd43073: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd43074: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd43075: begin  
rid<=0;
end
19'd43201: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=1;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=17971;
 end   
19'd43202: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=35;
   mapp<=70;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=20225;
 end   
19'd43203: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=93;
   mapp<=85;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=18090;
 end   
19'd43204: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=72;
   mapp<=52;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=14362;
 end   
19'd43205: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=16;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd43206: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=16;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd43207: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=28;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd43208: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=11;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd43209: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=25;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd43210: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd43211: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=88;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=38110;
 end   
19'd43212: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=21;
   mapp<=39;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=33871;
 end   
19'd43213: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=86;
   mapp<=44;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=36604;
 end   
19'd43214: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=8;
   mapp<=56;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=29749;
 end   
19'd43215: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=77;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd43216: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=28;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd43217: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=79;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd43218: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=47;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd43219: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=49;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd43220: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=80;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd43221: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd43363: begin  
rid<=1;
end
19'd43364: begin  
end
19'd43365: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd43366: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd43367: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd43368: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd43369: begin  
rid<=0;
end
19'd43501: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=19;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3180;
 end   
19'd43502: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=77;
   mapp<=26;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7150;
 end   
19'd43503: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=91;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6884;
 end   
19'd43504: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=47;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5154;
 end   
19'd43505: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=85;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd43506: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=84;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=6108;
 end   
19'd43507: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=54;
   mapp<=6;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=9238;
 end   
19'd43508: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=69;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=9077;
 end   
19'd43509: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=9;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=5769;
 end   
19'd43510: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=56;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd43511: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd43653: begin  
rid<=1;
end
19'd43654: begin  
end
19'd43655: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd43656: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd43657: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd43658: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd43659: begin  
rid<=0;
end
19'd43801: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=35;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13088;
 end   
19'd43802: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=90;
   mapp<=16;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10517;
 end   
19'd43803: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=77;
   mapp<=60;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=14451;
 end   
19'd43804: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=49;
   mapp<=97;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=16991;
 end   
19'd43805: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=5;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd43806: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=86;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd43807: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd43808: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=87;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=29882;
 end   
19'd43809: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=55;
   mapp<=43;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=22249;
 end   
19'd43810: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=82;
   mapp<=77;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=24500;
 end   
19'd43811: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=53;
   mapp<=30;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=27794;
 end   
19'd43812: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd43813: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=54;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd43814: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd43815: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd43957: begin  
rid<=1;
end
19'd43958: begin  
end
19'd43959: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd43960: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd43961: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd43962: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd43963: begin  
rid<=0;
end
19'd44101: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=54;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10367;
 end   
19'd44102: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=4;
   mapp<=10;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12618;
 end   
19'd44103: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=37;
   mapp<=40;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6760;
 end   
19'd44104: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=85;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd44105: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd44106: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd44107: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=51;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=18961;
 end   
19'd44108: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=29;
   mapp<=92;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20837;
 end   
19'd44109: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=37;
   mapp<=13;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=13544;
 end   
19'd44110: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=33;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd44111: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd44112: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd44113: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd44255: begin  
rid<=1;
end
19'd44256: begin  
end
19'd44257: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd44258: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd44259: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd44260: begin  
rid<=0;
end
19'd44401: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=68;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6214;
 end   
19'd44402: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=10;
   mapp<=57;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4716;
 end   
19'd44403: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=68;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6120;
 end   
19'd44404: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=8;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3031;
 end   
19'd44405: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=41;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5267;
 end   
19'd44406: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=32;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=4815;
 end   
19'd44407: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=37;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=7919;
 end   
19'd44408: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=84;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=12685;
 end   
19'd44409: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=99;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd44410: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=83;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=10161;
 end   
19'd44411: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=56;
   mapp<=69;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=11120;
 end   
19'd44412: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=92;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=8972;
 end   
19'd44413: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=40;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=9074;
 end   
19'd44414: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=87;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=6182;
 end   
19'd44415: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=12;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=5517;
 end   
19'd44416: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=10;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=9309;
 end   
19'd44417: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=20;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=15120;
 end   
19'd44418: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=35;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd44419: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd44561: begin  
rid<=1;
end
19'd44562: begin  
end
19'd44563: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd44564: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd44565: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd44566: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd44567: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd44568: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd44569: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd44570: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd44571: begin  
rid<=0;
end
19'd44701: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=34;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3298;
 end   
19'd44702: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2628;
 end   
19'd44703: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=74;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2536;
 end   
19'd44704: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=86;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7856;
 end   
19'd44705: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=33;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=5466;
 end   
19'd44706: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=78;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=9244;
 end   
19'd44707: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd44849: begin  
rid<=1;
end
19'd44850: begin  
end
19'd44851: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd44852: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd44853: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd44854: begin  
rid<=0;
end
19'd45001: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=4;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11334;
 end   
19'd45002: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=22;
   mapp<=49;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=19199;
 end   
19'd45003: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=55;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd45004: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=13;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd45005: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=62;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd45006: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=73;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd45007: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=84;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd45008: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=37;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=19637;
 end   
19'd45009: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=17;
   mapp<=22;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=33313;
 end   
19'd45010: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=6;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd45011: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=31;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd45012: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=97;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd45013: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=5;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd45014: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=36;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd45015: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd45157: begin  
rid<=1;
end
19'd45158: begin  
end
19'd45159: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd45160: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd45161: begin  
rid<=0;
end
19'd45301: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=96;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=26675;
 end   
19'd45302: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=55;
   mapp<=98;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=25050;
 end   
19'd45303: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=28;
   mapp<=85;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=23919;
 end   
19'd45304: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=38;
   mapp<=47;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=21493;
 end   
19'd45305: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=42;
   mapp<=84;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=21948;
 end   
19'd45306: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=28;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd45307: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=95;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd45308: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=42;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd45309: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd45310: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=6;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd45311: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=67;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd45312: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=65;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=41445;
 end   
19'd45313: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=39;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=36587;
 end   
19'd45314: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=6;
   mapp<=5;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=34921;
 end   
19'd45315: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=9;
   mapp<=46;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=38797;
 end   
19'd45316: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=92;
   mapp<=9;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=40711;
 end   
19'd45317: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=99;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd45318: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=75;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd45319: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=36;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd45320: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=61;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd45321: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=47;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd45322: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=18;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd45323: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd45465: begin  
rid<=1;
end
19'd45466: begin  
end
19'd45467: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd45468: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd45469: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd45470: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd45471: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd45472: begin  
rid<=0;
end
19'd45601: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=44;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=21869;
 end   
19'd45602: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=36;
   mapp<=96;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=23211;
 end   
19'd45603: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=37;
   mapp<=9;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=20539;
 end   
19'd45604: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=16;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd45605: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=93;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd45606: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=49;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd45607: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=71;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd45608: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=44;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd45609: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=77;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd45610: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd45611: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd45612: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=25;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=40224;
 end   
19'd45613: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=36;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=42005;
 end   
19'd45614: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=80;
   mapp<=90;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=36464;
 end   
19'd45615: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=16;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd45616: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=70;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd45617: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=84;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd45618: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=47;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd45619: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=28;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd45620: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=36;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd45621: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd45622: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd45623: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd45765: begin  
rid<=1;
end
19'd45766: begin  
end
19'd45767: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd45768: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd45769: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd45770: begin  
rid<=0;
end
19'd45901: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=64;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1472;
 end   
19'd45902: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=11;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=263;
 end   
19'd45903: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=40;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=940;
 end   
19'd45904: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=50;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1180;
 end   
19'd45905: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=4;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=132;
 end   
19'd45906: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=83;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=1959;
 end   
19'd45907: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=66;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=1578;
 end   
19'd45908: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=41;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=1013;
 end   
19'd45909: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=70;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=1690;
 end   
19'd45910: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=6;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=1742;
 end   
19'd45911: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=88;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=4223;
 end   
19'd45912: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=56;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=3460;
 end   
19'd45913: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=7;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=1495;
 end   
19'd45914: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=66;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=3102;
 end   
19'd45915: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=57;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=4524;
 end   
19'd45916: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=78;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=5088;
 end   
19'd45917: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=99;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=5468;
 end   
19'd45918: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=74;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=5020;
 end   
19'd45919: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd46061: begin  
rid<=1;
end
19'd46062: begin  
end
19'd46063: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd46064: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd46065: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd46066: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd46067: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd46068: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd46069: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd46070: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd46071: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd46072: begin  
rid<=0;
end
19'd46201: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=62;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5644;
 end   
19'd46202: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=2;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2110;
 end   
19'd46203: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=58;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3808;
 end   
19'd46204: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=96;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6016;
 end   
19'd46205: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=17;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1274;
 end   
19'd46206: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=90;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=5764;
 end   
19'd46207: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=67;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=4228;
 end   
19'd46208: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=7;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=572;
 end   
19'd46209: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=34;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=2280;
 end   
19'd46210: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd46211: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=79;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8751;
 end   
19'd46212: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=1;
   mapp<=26;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=4259;
 end   
19'd46213: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=95;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=11319;
 end   
19'd46214: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=6;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6504;
 end   
19'd46215: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=14;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=2430;
 end   
19'd46216: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=50;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=9800;
 end   
19'd46217: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=86;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=11101;
 end   
19'd46218: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=79;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=6889;
 end   
19'd46219: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=76;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=8306;
 end   
19'd46220: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd46221: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd46363: begin  
rid<=1;
end
19'd46364: begin  
end
19'd46365: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd46366: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd46367: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd46368: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd46369: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd46370: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd46371: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd46372: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd46373: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd46374: begin  
rid<=0;
end
19'd46501: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=61;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3904;
 end   
19'd46502: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=57;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3487;
 end   
19'd46503: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4290;
 end   
19'd46504: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=38;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=2348;
 end   
19'd46505: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=12;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=772;
 end   
19'd46506: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=44;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=2734;
 end   
19'd46507: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=39;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7024;
 end   
19'd46508: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=3487;
 end   
19'd46509: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=43;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=5967;
 end   
19'd46510: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=56;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=4532;
 end   
19'd46511: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=61;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=3151;
 end   
19'd46512: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=47;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=4567;
 end   
19'd46513: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd46655: begin  
rid<=1;
end
19'd46656: begin  
end
19'd46657: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd46658: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd46659: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd46660: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd46661: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd46662: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd46663: begin  
rid<=0;
end
19'd46801: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=13;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7747;
 end   
19'd46802: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=9;
   mapp<=79;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9427;
 end   
19'd46803: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=71;
   mapp<=18;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10630;
 end   
19'd46804: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=42;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd46805: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=39;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd46806: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=36;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd46807: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=21;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd46808: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd46809: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd46810: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=2;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=22178;
 end   
19'd46811: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=5;
   mapp<=34;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=19357;
 end   
19'd46812: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=38;
   mapp<=29;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=28861;
 end   
19'd46813: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=32;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd46814: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=65;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd46815: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=16;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd46816: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=81;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd46817: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd46818: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd46819: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd46961: begin  
rid<=1;
end
19'd46962: begin  
end
19'd46963: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd46964: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd46965: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd46966: begin  
rid<=0;
end
19'd47101: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=40;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4918;
 end   
19'd47102: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=16;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd47103: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=88;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd47104: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=19;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd47105: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=71;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=18030;
 end   
19'd47106: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=83;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd47107: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=64;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd47108: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=38;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd47109: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd47251: begin  
rid<=1;
end
19'd47252: begin  
end
19'd47253: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd47254: begin  
rid<=0;
end
19'd47401: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=16;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12915;
 end   
19'd47402: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=77;
   mapp<=1;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=14411;
 end   
19'd47403: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=52;
   mapp<=74;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=15792;
 end   
19'd47404: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=65;
   mapp<=33;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=18495;
 end   
19'd47405: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=91;
   mapp<=59;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=14345;
 end   
19'd47406: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=38;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd47407: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd47408: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd47409: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd47410: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd47411: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=34;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=29590;
 end   
19'd47412: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=68;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=30106;
 end   
19'd47413: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=41;
   mapp<=55;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=31832;
 end   
19'd47414: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=72;
   mapp<=87;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=33135;
 end   
19'd47415: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=68;
   mapp<=24;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=24768;
 end   
19'd47416: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=74;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd47417: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd47418: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd47419: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd47420: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd47421: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd47563: begin  
rid<=1;
end
19'd47564: begin  
end
19'd47565: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd47566: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd47567: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd47568: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd47569: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd47570: begin  
rid<=0;
end
19'd47701: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=15;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=495;
 end   
19'd47702: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=41;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=625;
 end   
19'd47703: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=45;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=695;
 end   
19'd47704: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=18;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=300;
 end   
19'd47705: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=24;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=2271;
 end   
19'd47706: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=52;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=1873;
 end   
19'd47707: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=46;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=1799;
 end   
19'd47708: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=56;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=1644;
 end   
19'd47709: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd47851: begin  
rid<=1;
end
19'd47852: begin  
end
19'd47853: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd47854: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd47855: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd47856: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd47857: begin  
rid<=0;
end
19'd48001: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=76;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6322;
 end   
19'd48002: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=27;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10746;
 end   
19'd48003: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=5;
   mapp<=34;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7990;
 end   
19'd48004: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=18;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd48005: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=91;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd48006: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=41;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd48007: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=11542;
 end   
19'd48008: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=17;
   mapp<=91;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=17776;
 end   
19'd48009: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=16;
   mapp<=71;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=18423;
 end   
19'd48010: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=43;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd48011: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=24;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd48012: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=64;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd48013: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd48155: begin  
rid<=1;
end
19'd48156: begin  
end
19'd48157: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd48158: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd48159: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd48160: begin  
rid<=0;
end
19'd48301: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=75;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3186;
 end   
19'd48302: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=46;
   mapp<=66;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2214;
 end   
19'd48303: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=32;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd48304: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=45;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7329;
 end   
19'd48305: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=3;
   mapp<=46;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=4873;
 end   
19'd48306: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=52;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd48307: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd48449: begin  
rid<=1;
end
19'd48450: begin  
end
19'd48451: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd48452: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd48453: begin  
rid<=0;
end
19'd48601: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=49;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6797;
 end   
19'd48602: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=50;
   mapp<=84;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3080;
 end   
19'd48603: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=5;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4149;
 end   
19'd48604: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=46;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4568;
 end   
19'd48605: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=25;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=7245;
 end   
19'd48606: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=70;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6784;
 end   
19'd48607: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=36;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=9948;
 end   
19'd48608: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=95;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=12917;
 end   
19'd48609: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=93;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=6941;
 end   
19'd48610: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=23;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=3997;
 end   
19'd48611: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=32;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd48612: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=10;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14653;
 end   
19'd48613: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=76;
   mapp<=96;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=16168;
 end   
19'd48614: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=92;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=14101;
 end   
19'd48615: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=50;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=16008;
 end   
19'd48616: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=90;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=21405;
 end   
19'd48617: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=95;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=17096;
 end   
19'd48618: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=52;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=17660;
 end   
19'd48619: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=50;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=17157;
 end   
19'd48620: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=15;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=11237;
 end   
19'd48621: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=36;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=11869;
 end   
19'd48622: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=61;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd48623: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd48765: begin  
rid<=1;
end
19'd48766: begin  
end
19'd48767: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd48768: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd48769: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd48770: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd48771: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd48772: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd48773: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd48774: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd48775: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd48776: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd48777: begin  
rid<=0;
end
19'd48901: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=66;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=20854;
 end   
19'd48902: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=16;
   mapp<=34;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=17190;
 end   
19'd48903: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=88;
   mapp<=50;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=14618;
 end   
19'd48904: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=25;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd48905: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=1;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd48906: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=10;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd48907: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=50;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd48908: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=82;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd48909: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd48910: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd48911: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=45;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=54733;
 end   
19'd48912: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=83;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=54481;
 end   
19'd48913: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=65;
   mapp<=38;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=45959;
 end   
19'd48914: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=96;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd48915: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=33;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd48916: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=90;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd48917: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=32;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd48918: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=89;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd48919: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd48920: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd48921: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd49063: begin  
rid<=1;
end
19'd49064: begin  
end
19'd49065: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd49066: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd49067: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd49068: begin  
rid<=0;
end
19'd49201: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=51;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11234;
 end   
19'd49202: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=18;
   mapp<=29;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7235;
 end   
19'd49203: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=63;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd49204: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=13;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd49205: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=7;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd49206: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=54;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd49207: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=76;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd49208: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=17;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd49209: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=11;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd49210: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=29;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd49211: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=58;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=40127;
 end   
19'd49212: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=64;
   mapp<=66;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=35652;
 end   
19'd49213: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=62;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd49214: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=10;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd49215: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=46;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd49216: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=65;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd49217: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=80;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd49218: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=65;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd49219: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=46;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd49220: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=40;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd49221: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd49363: begin  
rid<=1;
end
19'd49364: begin  
end
19'd49365: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd49366: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd49367: begin  
rid<=0;
end
19'd49501: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=6;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=572;
 end   
19'd49502: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=2;
   mapp<=94;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=742;
 end   
19'd49503: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=84;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=664;
 end   
19'd49504: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=70;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=480;
 end   
19'd49505: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=15;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=130;
 end   
19'd49506: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=62;
 end   
19'd49507: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd49508: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=54;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7340;
 end   
19'd49509: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=48;
   mapp<=33;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=3052;
 end   
19'd49510: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=11;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=4474;
 end   
19'd49511: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=67;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=4818;
 end   
19'd49512: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=15;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=3100;
 end   
19'd49513: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=45;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=6092;
 end   
19'd49514: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd49515: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd49657: begin  
rid<=1;
end
19'd49658: begin  
end
19'd49659: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd49660: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd49661: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd49662: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd49663: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd49664: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd49665: begin  
rid<=0;
end
19'd49801: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=9;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=792;
 end   
19'd49802: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=21;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=199;
 end   
19'd49803: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=92;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=848;
 end   
19'd49804: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=97;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=903;
 end   
19'd49805: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=97;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=913;
 end   
19'd49806: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=97;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5836;
 end   
19'd49807: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=71;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=7086;
 end   
19'd49808: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=58;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=6474;
 end   
19'd49809: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=22;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=3037;
 end   
19'd49810: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=59;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=6636;
 end   
19'd49811: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd49953: begin  
rid<=1;
end
19'd49954: begin  
end
19'd49955: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd49956: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd49957: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd49958: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd49959: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd49960: begin  
rid<=0;
end
19'd50101: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=8;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16782;
 end   
19'd50102: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=44;
   mapp<=20;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=13145;
 end   
19'd50103: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=69;
   mapp<=36;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=17042;
 end   
19'd50104: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=81;
   mapp<=84;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=18247;
 end   
19'd50105: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=79;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd50106: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=8;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd50107: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=7;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd50108: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=59;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd50109: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd50110: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd50111: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd50112: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=81;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=31576;
 end   
19'd50113: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=14;
   mapp<=49;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=29778;
 end   
19'd50114: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=49;
   mapp<=75;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=31321;
 end   
19'd50115: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=68;
   mapp<=26;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=33910;
 end   
19'd50116: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=38;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd50117: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=7;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd50118: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=93;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd50119: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=4;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd50120: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd50121: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd50122: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd50123: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd50265: begin  
rid<=1;
end
19'd50266: begin  
end
19'd50267: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd50268: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd50269: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd50270: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd50271: begin  
rid<=0;
end
19'd50401: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=79;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6997;
 end   
19'd50402: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=36;
   mapp<=55;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9285;
 end   
19'd50403: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=55;
   mapp<=41;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9823;
 end   
19'd50404: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=33;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd50405: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd50406: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd50407: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=70;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16445;
 end   
19'd50408: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=54;
   mapp<=30;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20485;
 end   
19'd50409: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=72;
   mapp<=52;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=26055;
 end   
19'd50410: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=76;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd50411: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd50412: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd50413: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd50555: begin  
rid<=1;
end
19'd50556: begin  
end
19'd50557: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd50558: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd50559: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd50560: begin  
rid<=0;
end
19'd50701: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=14;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=15972;
 end   
19'd50702: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=38;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd50703: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=57;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd50704: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=90;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd50705: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=38;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd50706: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=31;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=29906;
 end   
19'd50707: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=61;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd50708: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=19;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd50709: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=81;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd50710: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=90;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd50711: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd50853: begin  
rid<=1;
end
19'd50854: begin  
end
19'd50855: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd50856: begin  
rid<=0;
end
19'd51001: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=6;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4843;
 end   
19'd51002: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=22;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11994;
 end   
19'd51003: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=86;
   mapp<=2;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=15285;
 end   
19'd51004: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=94;
   mapp<=28;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=16971;
 end   
19'd51005: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=77;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd51006: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd51007: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd51008: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd51009: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=53;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=22039;
 end   
19'd51010: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=68;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=29688;
 end   
19'd51011: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=30;
   mapp<=47;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=28084;
 end   
19'd51012: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=55;
   mapp<=40;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=30498;
 end   
19'd51013: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=66;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd51014: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd51015: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd51016: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd51017: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd51159: begin  
rid<=1;
end
19'd51160: begin  
end
19'd51161: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd51162: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd51163: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd51164: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd51165: begin  
rid<=0;
end
19'd51301: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=23;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10526;
 end   
19'd51302: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=70;
   mapp<=18;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9470;
 end   
19'd51303: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=12;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd51304: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=50;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd51305: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=75;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd51306: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=11;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd51307: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=50;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd51308: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd51309: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=84;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=38949;
 end   
19'd51310: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=45;
   mapp<=88;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=35377;
 end   
19'd51311: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=87;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd51312: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=62;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd51313: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=43;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd51314: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=58;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd51315: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=59;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd51316: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd51317: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd51459: begin  
rid<=1;
end
19'd51460: begin  
end
19'd51461: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd51462: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd51463: begin  
rid<=0;
end
19'd51601: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=76;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10002;
 end   
19'd51602: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=16;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11232;
 end   
19'd51603: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=98;
   mapp<=41;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=13088;
 end   
19'd51604: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=83;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=9216;
 end   
19'd51605: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd51606: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd51607: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=75;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14773;
 end   
19'd51608: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=17;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=25981;
 end   
19'd51609: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=87;
   mapp<=5;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=19114;
 end   
19'd51610: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=97;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=23276;
 end   
19'd51611: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd51612: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd51613: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd51755: begin  
rid<=1;
end
19'd51756: begin  
end
19'd51757: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd51758: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd51759: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd51760: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd51761: begin  
rid<=0;
end
19'd51901: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=77;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13453;
 end   
19'd51902: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=86;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=16272;
 end   
19'd51903: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=81;
   mapp<=89;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=19631;
 end   
19'd51904: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=73;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=18444;
 end   
19'd51905: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd51906: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd51907: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=35;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=20933;
 end   
19'd51908: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=35;
   mapp<=22;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=25174;
 end   
19'd51909: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=83;
   mapp<=45;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=31026;
 end   
19'd51910: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=79;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=25263;
 end   
19'd51911: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd51912: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd51913: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd52055: begin  
rid<=1;
end
19'd52056: begin  
end
19'd52057: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd52058: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd52059: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd52060: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd52061: begin  
rid<=0;
end
19'd52201: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=36;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14566;
 end   
19'd52202: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=92;
   mapp<=85;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=13899;
 end   
19'd52203: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=65;
   mapp<=52;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=14120;
 end   
19'd52204: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=78;
   mapp<=21;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=14444;
 end   
19'd52205: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=60;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=18948;
 end   
19'd52206: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=82;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=13516;
 end   
19'd52207: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd52208: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd52209: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd52210: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=2;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=25052;
 end   
19'd52211: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=64;
   mapp<=96;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=25496;
 end   
19'd52212: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=39;
   mapp<=86;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=21344;
 end   
19'd52213: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=72;
   mapp<=11;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=22675;
 end   
19'd52214: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=76;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=23071;
 end   
19'd52215: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=47;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=18272;
 end   
19'd52216: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd52217: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd52218: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd52219: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd52361: begin  
rid<=1;
end
19'd52362: begin  
end
19'd52363: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd52364: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd52365: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd52366: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd52367: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd52368: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd52369: begin  
rid<=0;
end
19'd52501: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=80;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12261;
 end   
19'd52502: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=98;
   mapp<=54;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10424;
 end   
19'd52503: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=91;
   mapp<=59;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5670;
 end   
19'd52504: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=60;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7139;
 end   
19'd52505: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=10;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd52506: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=91;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd52507: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=36;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=23565;
 end   
19'd52508: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=99;
   mapp<=33;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=26282;
 end   
19'd52509: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=75;
   mapp<=75;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=19365;
 end   
19'd52510: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=90;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=19877;
 end   
19'd52511: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=76;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd52512: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=56;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd52513: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd52655: begin  
rid<=1;
end
19'd52656: begin  
end
19'd52657: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd52658: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd52659: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd52660: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd52661: begin  
rid<=0;
end
19'd52801: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=64;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11199;
 end   
19'd52802: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=85;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5573;
 end   
19'd52803: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=15;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4550;
 end   
19'd52804: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=42;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=10793;
 end   
19'd52805: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=95;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=11730;
 end   
19'd52806: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=66;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=9034;
 end   
19'd52807: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=56;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=10954;
 end   
19'd52808: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=86;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=8719;
 end   
19'd52809: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=37;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=10778;
 end   
19'd52810: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=98;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=8572;
 end   
19'd52811: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd52812: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=30;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=13541;
 end   
19'd52813: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=49;
   mapp<=8;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=7773;
 end   
19'd52814: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=40;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=8690;
 end   
19'd52815: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=60;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=13279;
 end   
19'd52816: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=14;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=14796;
 end   
19'd52817: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=54;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=11242;
 end   
19'd52818: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=12;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=13862;
 end   
19'd52819: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=52;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=12141;
 end   
19'd52820: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=38;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=12212;
 end   
19'd52821: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=6;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=9977;
 end   
19'd52822: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd52823: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd52965: begin  
rid<=1;
end
19'd52966: begin  
end
19'd52967: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd52968: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd52969: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd52970: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd52971: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd52972: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd52973: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd52974: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd52975: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd52976: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd52977: begin  
rid<=0;
end
19'd53101: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=21;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3530;
 end   
19'd53102: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=45;
   mapp<=38;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5226;
 end   
19'd53103: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=91;
   mapp<=17;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4488;
 end   
19'd53104: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=69;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=2545;
 end   
19'd53105: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=39;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1956;
 end   
19'd53106: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=8;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=3678;
 end   
19'd53107: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=65;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=4502;
 end   
19'd53108: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=62;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=5027;
 end   
19'd53109: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=73;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=5297;
 end   
19'd53110: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=81;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd53111: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd53112: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=8;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=4933;
 end   
19'd53113: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=15;
   mapp<=53;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=7996;
 end   
19'd53114: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=29;
   mapp<=8;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=10061;
 end   
19'd53115: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=66;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=10868;
 end   
19'd53116: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=89;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=10046;
 end   
19'd53117: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=63;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=10730;
 end   
19'd53118: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=71;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=10484;
 end   
19'd53119: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=41;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=10329;
 end   
19'd53120: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=59;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=10289;
 end   
19'd53121: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=31;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd53122: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=72;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd53123: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd53265: begin  
rid<=1;
end
19'd53266: begin  
end
19'd53267: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd53268: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd53269: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd53270: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd53271: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd53272: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd53273: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd53274: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd53275: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd53276: begin  
rid<=0;
end
19'd53401: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=36;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16698;
 end   
19'd53402: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=78;
   mapp<=70;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=16420;
 end   
19'd53403: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=6;
   mapp<=68;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=14066;
 end   
19'd53404: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=27;
   mapp<=99;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=19728;
 end   
19'd53405: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=13;
   mapp<=55;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=20572;
 end   
19'd53406: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=23;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd53407: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=71;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd53408: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=27;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd53409: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=73;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd53410: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=61;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd53411: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=73;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd53412: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=95;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=29018;
 end   
19'd53413: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=95;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=27866;
 end   
19'd53414: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=13;
   mapp<=87;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=27874;
 end   
19'd53415: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=6;
   mapp<=17;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=33685;
 end   
19'd53416: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=70;
   mapp<=63;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=29787;
 end   
19'd53417: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=59;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd53418: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=5;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd53419: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=96;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd53420: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=33;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd53421: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd53422: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=52;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd53423: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd53565: begin  
rid<=1;
end
19'd53566: begin  
end
19'd53567: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd53568: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd53569: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd53570: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd53571: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd53572: begin  
rid<=0;
end
19'd53701: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=44;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=20514;
 end   
19'd53702: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=7;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=21974;
 end   
19'd53703: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=71;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd53704: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=87;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd53705: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=99;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd53706: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=19;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd53707: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=57;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=40206;
 end   
19'd53708: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=90;
   mapp<=15;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=42852;
 end   
19'd53709: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=59;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd53710: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=57;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd53711: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=86;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd53712: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=9;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd53713: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd53855: begin  
rid<=1;
end
19'd53856: begin  
end
19'd53857: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd53858: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd53859: begin  
rid<=0;
end
19'd54001: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=35;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2317;
 end   
19'd54002: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=28;
   mapp<=59;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2439;
 end   
19'd54003: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd54004: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=56;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=4481;
 end   
19'd54005: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=31;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8386;
 end   
19'd54006: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd54007: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd54149: begin  
rid<=1;
end
19'd54150: begin  
end
19'd54151: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd54152: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd54153: begin  
rid<=0;
end
19'd54301: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=74;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=18014;
 end   
19'd54302: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=38;
   mapp<=43;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9769;
 end   
19'd54303: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=83;
   mapp<=74;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=16809;
 end   
19'd54304: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=58;
   mapp<=16;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=10059;
 end   
19'd54305: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=95;
   mapp<=24;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=17310;
 end   
19'd54306: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=11;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=15453;
 end   
19'd54307: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=85;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=25410;
 end   
19'd54308: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd54309: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd54310: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd54311: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd54312: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=58;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=23374;
 end   
19'd54313: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=18;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=17264;
 end   
19'd54314: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=57;
   mapp<=31;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=22285;
 end   
19'd54315: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=61;
   mapp<=3;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=17899;
 end   
19'd54316: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=20;
   mapp<=32;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=29336;
 end   
19'd54317: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=22221;
 end   
19'd54318: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=90;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=32871;
 end   
19'd54319: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd54320: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd54321: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd54322: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd54323: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd54465: begin  
rid<=1;
end
19'd54466: begin  
end
19'd54467: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd54468: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd54469: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd54470: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd54471: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd54472: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd54473: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd54474: begin  
rid<=0;
end
19'd54601: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=92;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3820;
 end   
19'd54602: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=82;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3220;
 end   
19'd54603: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=67;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1531;
 end   
19'd54604: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=20;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=2146;
 end   
19'd54605: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=58;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3162;
 end   
19'd54606: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=74;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=3796;
 end   
19'd54607: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=87;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd54608: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=64;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=15148;
 end   
19'd54609: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=64;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=10398;
 end   
19'd54610: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=14;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=6665;
 end   
19'd54611: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=46;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=13940;
 end   
19'd54612: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=90;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=13697;
 end   
19'd54613: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=25;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=10711;
 end   
19'd54614: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=55;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd54615: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd54757: begin  
rid<=1;
end
19'd54758: begin  
end
19'd54759: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd54760: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd54761: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd54762: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd54763: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd54764: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd54765: begin  
rid<=0;
end
19'd54901: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=79;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=21555;
 end   
19'd54902: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=91;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd54903: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=66;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd54904: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=87;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd54905: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=8;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd54906: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=26;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd54907: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=25;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd54908: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=59;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd54909: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=60;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=38402;
 end   
19'd54910: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=51;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd54911: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=8;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd54912: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=78;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd54913: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=94;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd54914: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=89;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd54915: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=24;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd54916: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=76;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd54917: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd55059: begin  
rid<=1;
end
19'd55060: begin  
end
19'd55061: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd55062: begin  
rid<=0;
end
19'd55201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=2;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3822;
 end   
19'd55202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=44;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6332;
 end   
19'd55203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=23;
   mapp<=19;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5073;
 end   
19'd55204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=39;
   mapp<=1;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4699;
 end   
19'd55205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=9;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3574;
 end   
19'd55206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=27;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6767;
 end   
19'd55207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=37;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=9876;
 end   
19'd55208: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=86;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd55209: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd55210: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=27;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd55211: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=15;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=10399;
 end   
19'd55212: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=44;
   mapp<=23;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18119;
 end   
19'd55213: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=36;
   mapp<=99;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=17930;
 end   
19'd55214: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=69;
   mapp<=14;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=19590;
 end   
19'd55215: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=78;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=17174;
 end   
19'd55216: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=76;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=19137;
 end   
19'd55217: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=58;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=20146;
 end   
19'd55218: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=52;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd55219: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=46;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd55220: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd55221: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd55363: begin  
rid<=1;
end
19'd55364: begin  
end
19'd55365: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd55366: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd55367: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd55368: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd55369: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd55370: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd55371: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd55372: begin  
rid<=0;
end
19'd55501: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=16;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=21438;
 end   
19'd55502: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=24;
   mapp<=88;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=27633;
 end   
19'd55503: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=29;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd55504: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=42;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd55505: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=84;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd55506: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=72;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd55507: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=49;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd55508: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=96;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd55509: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=26;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd55510: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=82;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd55511: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=54;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=36757;
 end   
19'd55512: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=43;
   mapp<=75;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=40668;
 end   
19'd55513: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=24;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd55514: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=99;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd55515: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=22;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd55516: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=21;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd55517: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=33;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd55518: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=13;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd55519: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=17;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd55520: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=93;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd55521: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd55663: begin  
rid<=1;
end
19'd55664: begin  
end
19'd55665: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd55666: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd55667: begin  
rid<=0;
end
19'd55801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=95;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12776;
 end   
19'd55802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=26;
   mapp<=74;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11976;
 end   
19'd55803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=20;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd55804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=91;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd55805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=88;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd55806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd55807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=22;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=23247;
 end   
19'd55808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=76;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=23143;
 end   
19'd55809: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=37;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd55810: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=16;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd55811: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=3;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd55812: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd55813: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd55955: begin  
rid<=1;
end
19'd55956: begin  
end
19'd55957: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd55958: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd55959: begin  
rid<=0;
end
19'd56101: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=22;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9053;
 end   
19'd56102: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=2;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd56103: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=2;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd56104: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=69;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd56105: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=74;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17237;
 end   
19'd56106: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=26;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd56107: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=63;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd56108: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=34;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd56109: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd56251: begin  
rid<=1;
end
19'd56252: begin  
end
19'd56253: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd56254: begin  
rid<=0;
end
19'd56401: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=37;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5349;
 end   
19'd56402: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=95;
   mapp<=3;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8448;
 end   
19'd56403: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=79;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd56404: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=61;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd56405: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=44;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd56406: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=59;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd56407: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=92;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=21000;
 end   
19'd56408: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=72;
   mapp<=7;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=22699;
 end   
19'd56409: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=28;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd56410: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=96;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd56411: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=11;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd56412: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=35;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd56413: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd56555: begin  
rid<=1;
end
19'd56556: begin  
end
19'd56557: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd56558: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd56559: begin  
rid<=0;
end
19'd56701: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=24;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14899;
 end   
19'd56702: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=20;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=18733;
 end   
19'd56703: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=26;
   mapp<=56;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=21780;
 end   
19'd56704: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=6;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd56705: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=83;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd56706: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=45;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd56707: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=74;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd56708: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=91;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd56709: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd56710: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=23;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=23478;
 end   
19'd56711: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=52;
   mapp<=64;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=29057;
 end   
19'd56712: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=25;
   mapp<=4;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=29877;
 end   
19'd56713: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=11;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd56714: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=42;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd56715: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=24;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd56716: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=49;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd56717: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=35;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd56718: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=90;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd56719: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd56861: begin  
rid<=1;
end
19'd56862: begin  
end
19'd56863: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd56864: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd56865: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd56866: begin  
rid<=0;
end
19'd57001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=79;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7756;
 end   
19'd57002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=2;
   mapp<=4;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1155;
 end   
19'd57003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=83;
   mapp<=41;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10000;
 end   
19'd57004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd57005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd57006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=47;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=13320;
 end   
19'd57007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=5;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=11629;
 end   
19'd57008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=90;
   mapp<=12;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=16549;
 end   
19'd57009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd57010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd57011: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd57153: begin  
rid<=1;
end
19'd57154: begin  
end
19'd57155: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd57156: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd57157: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd57158: begin  
rid<=0;
end
19'd57301: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=80;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7193;
 end   
19'd57302: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=71;
   mapp<=39;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6160;
 end   
19'd57303: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=78;
   mapp<=28;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5332;
 end   
19'd57304: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=40;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4678;
 end   
19'd57305: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=56;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4712;
 end   
19'd57306: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=48;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd57307: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=44;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd57308: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=98;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12803;
 end   
19'd57309: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=16;
   mapp<=25;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=9030;
 end   
19'd57310: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=80;
   mapp<=10;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=9947;
 end   
19'd57311: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=15;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=7213;
 end   
19'd57312: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=64;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=8962;
 end   
19'd57313: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=26;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd57314: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=72;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd57315: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd57457: begin  
rid<=1;
end
19'd57458: begin  
end
19'd57459: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd57460: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd57461: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd57462: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd57463: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd57464: begin  
rid<=0;
end
19'd57601: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=36;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3117;
 end   
19'd57602: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=33;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2741;
 end   
19'd57603: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=5;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd57604: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=38;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8503;
 end   
19'd57605: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=65;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=10444;
 end   
19'd57606: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=64;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd57607: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd57749: begin  
rid<=1;
end
19'd57750: begin  
end
19'd57751: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd57752: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd57753: begin  
rid<=0;
end
19'd57901: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=62;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=17289;
 end   
19'd57902: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=69;
   mapp<=8;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=18089;
 end   
19'd57903: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=49;
   mapp<=96;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=22504;
 end   
19'd57904: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=18;
   mapp<=38;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=20287;
 end   
19'd57905: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=67;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd57906: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=58;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd57907: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=43;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd57908: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd57909: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd57910: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd57911: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=47;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=30810;
 end   
19'd57912: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=96;
   mapp<=3;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=33729;
 end   
19'd57913: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=66;
   mapp<=90;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=37056;
 end   
19'd57914: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=30;
   mapp<=86;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=30679;
 end   
19'd57915: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=65;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd57916: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=52;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd57917: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd57918: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd57919: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd57920: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd57921: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd58063: begin  
rid<=1;
end
19'd58064: begin  
end
19'd58065: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd58066: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd58067: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd58068: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd58069: begin  
rid<=0;
end
19'd58201: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=12;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3344;
 end   
19'd58202: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=34;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4124;
 end   
19'd58203: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=97;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3870;
 end   
19'd58204: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=79;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1794;
 end   
19'd58205: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=24;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1280;
 end   
19'd58206: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=28;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=2426;
 end   
19'd58207: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=60;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=2752;
 end   
19'd58208: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=58;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=1616;
 end   
19'd58209: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=25;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=2658;
 end   
19'd58210: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd58211: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=60;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=9569;
 end   
19'd58212: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=45;
   mapp<=69;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=11054;
 end   
19'd58213: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=62;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=10740;
 end   
19'd58214: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=70;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6489;
 end   
19'd58215: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=11;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=3515;
 end   
19'd58216: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=35;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=8576;
 end   
19'd58217: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=90;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=8647;
 end   
19'd58218: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=11;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=5156;
 end   
19'd58219: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=64;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=8748;
 end   
19'd58220: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd58221: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd58363: begin  
rid<=1;
end
19'd58364: begin  
end
19'd58365: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd58366: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd58367: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd58368: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd58369: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd58370: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd58371: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd58372: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd58373: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd58374: begin  
rid<=0;
end
19'd58501: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=15;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=21099;
 end   
19'd58502: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=79;
   mapp<=17;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=25888;
 end   
19'd58503: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=37;
   mapp<=65;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=16129;
 end   
19'd58504: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=88;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd58505: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=69;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd58506: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=86;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd58507: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=30;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd58508: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=9;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd58509: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=11;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=34706;
 end   
19'd58510: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=54;
   mapp<=21;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=39508;
 end   
19'd58511: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=93;
   mapp<=19;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=32231;
 end   
19'd58512: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=84;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd58513: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=57;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd58514: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=99;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd58515: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=36;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd58516: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=29;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd58517: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd58659: begin  
rid<=1;
end
19'd58660: begin  
end
19'd58661: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd58662: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd58663: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd58664: begin  
rid<=0;
end
19'd58801: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=17;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=26513;
 end   
19'd58802: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=77;
   mapp<=65;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=20859;
 end   
19'd58803: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=60;
   mapp<=34;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=17952;
 end   
19'd58804: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=5;
   mapp<=49;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=21359;
 end   
19'd58805: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=53;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd58806: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=91;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd58807: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=62;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd58808: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=76;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd58809: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd58810: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd58811: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd58812: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=44;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=44216;
 end   
19'd58813: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=59;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=39336;
 end   
19'd58814: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=66;
   mapp<=34;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=36045;
 end   
19'd58815: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=85;
   mapp<=16;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=42145;
 end   
19'd58816: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=39;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd58817: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=18;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd58818: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=7;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd58819: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=68;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd58820: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd58821: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd58822: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd58823: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd58965: begin  
rid<=1;
end
19'd58966: begin  
end
19'd58967: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd58968: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd58969: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd58970: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd58971: begin  
rid<=0;
end
19'd59101: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=20;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4105;
 end   
19'd59102: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=35;
   mapp<=99;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10832;
 end   
19'd59103: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=98;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12264;
 end   
19'd59104: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=92;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4558;
 end   
19'd59105: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=16;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=8670;
 end   
19'd59106: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=82;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=5545;
 end   
19'd59107: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=29;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=2572;
 end   
19'd59108: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd59109: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=83;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14744;
 end   
19'd59110: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=99;
   mapp<=58;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18703;
 end   
19'd59111: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=35;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=17635;
 end   
19'd59112: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=57;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=11981;
 end   
19'd59113: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=70;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=16918;
 end   
19'd59114: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=71;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=12170;
 end   
19'd59115: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=42;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=9690;
 end   
19'd59116: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=80;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd59117: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd59259: begin  
rid<=1;
end
19'd59260: begin  
end
19'd59261: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd59262: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd59263: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd59264: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd59265: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd59266: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd59267: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd59268: begin  
rid<=0;
end
19'd59401: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=28;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9548;
 end   
19'd59402: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=78;
   mapp<=86;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5772;
 end   
19'd59403: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=60;
   mapp<=3;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5240;
 end   
19'd59404: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=52;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4990;
 end   
19'd59405: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=18;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=8374;
 end   
19'd59406: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd59407: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd59408: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=41;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17403;
 end   
19'd59409: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=38;
   mapp<=49;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18118;
 end   
19'd59410: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=93;
   mapp<=64;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=13512;
 end   
19'd59411: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=85;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=14764;
 end   
19'd59412: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=26;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=15047;
 end   
19'd59413: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd59414: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd59415: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd59557: begin  
rid<=1;
end
19'd59558: begin  
end
19'd59559: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd59560: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd59561: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd59562: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd59563: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd59564: begin  
rid<=0;
end
19'd59701: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=35;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10875;
 end   
19'd59702: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=9;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd59703: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=96;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd59704: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=84;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=22943;
 end   
19'd59705: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=23;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd59706: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=99;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd59707: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd59849: begin  
rid<=1;
end
19'd59850: begin  
end
19'd59851: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd59852: begin  
rid<=0;
end
19'd60001: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=6;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=252;
 end   
19'd60002: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=50;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2110;
 end   
19'd60003: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=87;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3674;
 end   
19'd60004: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=69;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=3012;
 end   
19'd60005: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=23;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=3030;
 end   
19'd60006: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=88;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=7194;
 end   
19'd60007: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd60149: begin  
rid<=1;
end
19'd60150: begin  
end
19'd60151: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd60152: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd60153: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd60154: begin  
rid<=0;
end
19'd60301: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=58;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=0;
 end   
19'd60302: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=6;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10;
 end   
19'd60303: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=38;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=20;
 end   
19'd60304: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=63;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=30;
 end   
19'd60305: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=20;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=40;
 end   
19'd60306: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=66;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=50;
 end   
19'd60307: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=85;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=4930;
 end   
19'd60308: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=23;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=1344;
 end   
19'd60309: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=29;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=1702;
 end   
19'd60310: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=98;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=5714;
 end   
19'd60311: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=56;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=3288;
 end   
19'd60312: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=70;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=4110;
 end   
19'd60313: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd60455: begin  
rid<=1;
end
19'd60456: begin  
end
19'd60457: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd60458: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd60459: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd60460: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd60461: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd60462: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd60463: begin  
rid<=0;
end
19'd60601: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=45;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=31074;
 end   
19'd60602: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=54;
   mapp<=88;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=28509;
 end   
19'd60603: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=58;
   mapp<=19;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=26414;
 end   
19'd60604: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=58;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd60605: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=94;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd60606: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=91;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd60607: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=41;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd60608: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=37;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd60609: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd60610: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd60611: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=53;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=56427;
 end   
19'd60612: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=27;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=51013;
 end   
19'd60613: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=85;
   mapp<=75;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=51692;
 end   
19'd60614: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=26;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd60615: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=70;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd60616: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=36;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd60617: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=81;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd60618: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=70;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd60619: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd60620: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd60621: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd60763: begin  
rid<=1;
end
19'd60764: begin  
end
19'd60765: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd60766: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd60767: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd60768: begin  
rid<=0;
end
19'd60901: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=51;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12627;
 end   
19'd60902: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=31;
   mapp<=99;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=13230;
 end   
19'd60903: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=17;
   mapp<=35;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=13702;
 end   
19'd60904: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=33;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd60905: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=71;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd60906: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=76;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd60907: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=29;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd60908: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=28;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=22260;
 end   
19'd60909: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=16;
   mapp<=44;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=23199;
 end   
19'd60910: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=34;
   mapp<=42;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=24186;
 end   
19'd60911: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=99;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd60912: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=57;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd60913: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=40;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd60914: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=81;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd60915: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd61057: begin  
rid<=1;
end
19'd61058: begin  
end
19'd61059: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd61060: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd61061: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd61062: begin  
rid<=0;
end
19'd61201: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=63;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5172;
 end   
19'd61202: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=45;
   mapp<=49;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7426;
 end   
19'd61203: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=26;
   mapp<=39;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8882;
 end   
19'd61204: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=99;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=12216;
 end   
19'd61205: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd61206: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd61207: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=95;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12157;
 end   
19'd61208: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=45;
   mapp<=24;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=19671;
 end   
19'd61209: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=70;
   mapp<=83;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=23222;
 end   
19'd61210: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=89;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=23926;
 end   
19'd61211: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd61212: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd61213: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd61355: begin  
rid<=1;
end
19'd61356: begin  
end
19'd61357: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd61358: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd61359: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd61360: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd61361: begin  
rid<=0;
end
19'd61501: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=65;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=17816;
 end   
19'd61502: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=14;
   mapp<=52;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=17741;
 end   
19'd61503: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=80;
   mapp<=24;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=15290;
 end   
19'd61504: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=58;
   mapp<=73;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=19627;
 end   
19'd61505: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=58;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd61506: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=24;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd61507: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=8;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd61508: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=11;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd61509: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd61510: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd61511: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd61512: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=75;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=39009;
 end   
19'd61513: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=84;
   mapp<=17;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=39349;
 end   
19'd61514: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=82;
   mapp<=28;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=41016;
 end   
19'd61515: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=11;
   mapp<=90;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=45043;
 end   
19'd61516: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=6;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd61517: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=68;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd61518: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=44;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd61519: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=26;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd61520: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd61521: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd61522: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd61523: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd61665: begin  
rid<=1;
end
19'd61666: begin  
end
19'd61667: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd61668: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd61669: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd61670: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd61671: begin  
rid<=0;
end
19'd61801: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=65;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8822;
 end   
19'd61802: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=12;
   mapp<=88;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6998;
 end   
19'd61803: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=47;
   mapp<=38;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10634;
 end   
19'd61804: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=46;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=11430;
 end   
19'd61805: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=59;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=12742;
 end   
19'd61806: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=52;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=13210;
 end   
19'd61807: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=71;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=11900;
 end   
19'd61808: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=56;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd61809: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=10;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd61810: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=70;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17032;
 end   
19'd61811: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=45;
   mapp<=66;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=13613;
 end   
19'd61812: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=25;
   mapp<=50;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=18927;
 end   
19'd61813: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=48;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=22750;
 end   
19'd61814: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=74;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=23994;
 end   
19'd61815: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=74;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=21716;
 end   
19'd61816: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=43;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=18065;
 end   
19'd61817: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=29;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd61818: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=36;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd61819: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd61961: begin  
rid<=1;
end
19'd61962: begin  
end
19'd61963: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd61964: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd61965: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd61966: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd61967: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd61968: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd61969: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd61970: begin  
rid<=0;
end
19'd62101: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=24;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14928;
 end   
19'd62102: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=34;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=13040;
 end   
19'd62103: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=75;
   mapp<=1;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=16532;
 end   
19'd62104: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=37;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd62105: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=76;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd62106: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd62107: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=24;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd62108: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=64;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd62109: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd62110: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd62111: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=71;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=46905;
 end   
19'd62112: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=90;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=43916;
 end   
19'd62113: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=84;
   mapp<=25;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=39352;
 end   
19'd62114: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=19;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd62115: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=79;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd62116: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=95;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd62117: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=58;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd62118: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=7;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd62119: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd62120: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd62121: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd62263: begin  
rid<=1;
end
19'd62264: begin  
end
19'd62265: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd62266: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd62267: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd62268: begin  
rid<=0;
end
19'd62401: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=89;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=19554;
 end   
19'd62402: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=25;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=22039;
 end   
19'd62403: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=29;
   mapp<=20;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=20408;
 end   
19'd62404: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=28;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd62405: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=39;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd62406: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=27;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd62407: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=94;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd62408: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=90;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd62409: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd62410: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd62411: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=43;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=40661;
 end   
19'd62412: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=39;
   mapp<=54;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=39882;
 end   
19'd62413: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=1;
   mapp<=17;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=42667;
 end   
19'd62414: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=93;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd62415: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=27;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd62416: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=69;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd62417: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=93;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd62418: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=33;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd62419: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd62420: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd62421: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd62563: begin  
rid<=1;
end
19'd62564: begin  
end
19'd62565: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd62566: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd62567: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd62568: begin  
rid<=0;
end
19'd62701: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=17;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7554;
 end   
19'd62702: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=7;
   mapp<=26;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=13283;
 end   
19'd62703: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=20;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd62704: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=45;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd62705: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=66;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd62706: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=21;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd62707: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=82;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd62708: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=43;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=26499;
 end   
19'd62709: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=63;
   mapp<=6;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=31092;
 end   
19'd62710: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=71;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd62711: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=92;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd62712: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=35;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd62713: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=17;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd62714: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd62715: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd62857: begin  
rid<=1;
end
19'd62858: begin  
end
19'd62859: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd62860: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd62861: begin  
rid<=0;
end
19'd63001: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=53;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6981;
 end   
19'd63002: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=51;
   mapp<=52;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7750;
 end   
19'd63003: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=94;
   mapp<=22;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6623;
 end   
19'd63004: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=41;
   mapp<=28;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6754;
 end   
19'd63005: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=30;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=9424;
 end   
19'd63006: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd63007: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd63008: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd63009: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=58;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14075;
 end   
19'd63010: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=2;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=19248;
 end   
19'd63011: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=53;
   mapp<=20;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=16308;
 end   
19'd63012: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=49;
   mapp<=44;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=14200;
 end   
19'd63013: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=88;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=15469;
 end   
19'd63014: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd63015: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd63016: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd63017: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd63159: begin  
rid<=1;
end
19'd63160: begin  
end
19'd63161: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd63162: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd63163: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd63164: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd63165: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd63166: begin  
rid<=0;
end
19'd63301: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=26;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9511;
 end   
19'd63302: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=30;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd63303: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=9;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd63304: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=20;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd63305: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=35;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd63306: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=43;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd63307: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=31;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd63308: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=74;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd63309: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=2;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd63310: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd63311: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=54;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=36310;
 end   
19'd63312: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=82;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd63313: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=33;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd63314: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=88;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd63315: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=55;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd63316: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=60;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd63317: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=45;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd63318: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=23;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd63319: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=42;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd63320: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=59;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd63321: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd63463: begin  
rid<=1;
end
19'd63464: begin  
end
19'd63465: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd63466: begin  
rid<=0;
end
19'd63601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=79;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9538;
 end   
19'd63602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=7;
   mapp<=84;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=13433;
 end   
19'd63603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=13;
   mapp<=89;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=14551;
 end   
19'd63604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=60;
   mapp<=68;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=12092;
 end   
19'd63605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd63606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd63607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd63608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=36;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=24363;
 end   
19'd63609: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=53;
   mapp<=46;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=26742;
 end   
19'd63610: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=49;
   mapp<=71;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=27305;
 end   
19'd63611: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=88;
   mapp<=82;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=23658;
 end   
19'd63612: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd63613: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd63614: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd63615: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd63757: begin  
rid<=1;
end
19'd63758: begin  
end
19'd63759: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd63760: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd63761: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd63762: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd63763: begin  
rid<=0;
end
19'd63901: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=85;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4335;
 end   
19'd63902: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=90;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7660;
 end   
19'd63903: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=39;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3335;
 end   
19'd63904: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=46;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3940;
 end   
19'd63905: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=62;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5310;
 end   
19'd63906: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=75;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6425;
 end   
19'd63907: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=24;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=2100;
 end   
19'd63908: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=78;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=6700;
 end   
19'd63909: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=29;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=4422;
 end   
19'd63910: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=81;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=10009;
 end   
19'd63911: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=77;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=5568;
 end   
19'd63912: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=50;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=5390;
 end   
19'd63913: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=48;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=6702;
 end   
19'd63914: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=70;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=8455;
 end   
19'd63915: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=94;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=4826;
 end   
19'd63916: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=16;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=7164;
 end   
19'd63917: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd64059: begin  
rid<=1;
end
19'd64060: begin  
end
19'd64061: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd64062: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd64063: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd64064: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd64065: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd64066: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd64067: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd64068: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd64069: begin  
rid<=0;
end
19'd64201: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=67;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1005;
 end   
19'd64202: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4834;
 end   
19'd64203: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=52;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3504;
 end   
19'd64204: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=62;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4184;
 end   
19'd64205: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=21;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1447;
 end   
19'd64206: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=89;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=3497;
 end   
19'd64207: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=65;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=10619;
 end   
19'd64208: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=29;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=6085;
 end   
19'd64209: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=59;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=9435;
 end   
19'd64210: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=82;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=8745;
 end   
19'd64211: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd64353: begin  
rid<=1;
end
19'd64354: begin  
end
19'd64355: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd64356: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd64357: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd64358: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd64359: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd64360: begin  
rid<=0;
end
19'd64501: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=3;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8881;
 end   
19'd64502: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=61;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7228;
 end   
19'd64503: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=96;
   mapp<=66;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10330;
 end   
19'd64504: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=32;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7423;
 end   
19'd64505: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd64506: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd64507: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=13;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14104;
 end   
19'd64508: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=65;
   mapp<=50;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=13198;
 end   
19'd64509: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=45;
   mapp<=32;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=18171;
 end   
19'd64510: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=72;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=15474;
 end   
19'd64511: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd64512: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd64513: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd64655: begin  
rid<=1;
end
19'd64656: begin  
end
19'd64657: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd64658: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd64659: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd64660: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd64661: begin  
rid<=0;
end
19'd64801: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=96;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3262;
 end   
19'd64802: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=4;
   mapp<=70;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3181;
 end   
19'd64803: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=14;
   mapp<=21;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7552;
 end   
19'd64804: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=99;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4951;
 end   
19'd64805: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=10;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6242;
 end   
19'd64806: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=69;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd64807: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=52;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd64808: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=30;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12818;
 end   
19'd64809: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=82;
   mapp<=71;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=14562;
 end   
19'd64810: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=61;
   mapp<=44;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=18676;
 end   
19'd64811: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=95;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=14801;
 end   
19'd64812: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=51;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=16365;
 end   
19'd64813: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=66;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd64814: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=83;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd64815: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd64957: begin  
rid<=1;
end
19'd64958: begin  
end
19'd64959: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd64960: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd64961: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd64962: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd64963: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd64964: begin  
rid<=0;
end
19'd65101: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=95;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6840;
 end   
19'd65102: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=6;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=442;
 end   
19'd65103: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=14;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1028;
 end   
19'd65104: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=52;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3774;
 end   
19'd65105: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=84;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6088;
 end   
19'd65106: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=5;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=410;
 end   
19'd65107: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=12;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=924;
 end   
19'd65108: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=41;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7701;
 end   
19'd65109: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=75;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=2017;
 end   
19'd65110: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=90;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=2918;
 end   
19'd65111: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=25;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=4299;
 end   
19'd65112: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=11;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=6319;
 end   
19'd65113: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=67;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=1817;
 end   
19'd65114: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=82;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=2646;
 end   
19'd65115: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd65257: begin  
rid<=1;
end
19'd65258: begin  
end
19'd65259: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd65260: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd65261: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd65262: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd65263: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd65264: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd65265: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd65266: begin  
rid<=0;
end
19'd65401: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=5;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1015;
 end   
19'd65402: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=11;
   mapp<=50;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1129;
 end   
19'd65403: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=79;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1163;
 end   
19'd65404: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=68;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1184;
 end   
19'd65405: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=74;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1334;
 end   
19'd65406: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=84;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=789;
 end   
19'd65407: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=29;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=590;
 end   
19'd65408: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=35;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=905;
 end   
19'd65409: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd65410: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=67;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7179;
 end   
19'd65411: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=24;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=2737;
 end   
19'd65412: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=50;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=4513;
 end   
19'd65413: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=16;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=2256;
 end   
19'd65414: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=60;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=5354;
 end   
19'd65415: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=1;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=856;
 end   
19'd65416: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=59;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=4543;
 end   
19'd65417: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=9;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=1508;
 end   
19'd65418: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd65419: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd65561: begin  
rid<=1;
end
19'd65562: begin  
end
19'd65563: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd65564: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd65565: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd65566: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd65567: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd65568: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd65569: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd65570: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd65571: begin  
rid<=0;
end
19'd65701: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=48;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1920;
 end   
19'd65702: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=55;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2210;
 end   
19'd65703: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=7;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=300;
 end   
19'd65704: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=49;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1990;
 end   
19'd65705: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=91;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3680;
 end   
19'd65706: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=60;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=2450;
 end   
19'd65707: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=82;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=3340;
 end   
19'd65708: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=19;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=2604;
 end   
19'd65709: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=70;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=4730;
 end   
19'd65710: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=79;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=3144;
 end   
19'd65711: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=25;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=2890;
 end   
19'd65712: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=19;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=4364;
 end   
19'd65713: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=9;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=2774;
 end   
19'd65714: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=1;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=3376;
 end   
19'd65715: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd65857: begin  
rid<=1;
end
19'd65858: begin  
end
19'd65859: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd65860: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd65861: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd65862: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd65863: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd65864: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd65865: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd65866: begin  
rid<=0;
end
19'd66001: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=70;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=19085;
 end   
19'd66002: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=51;
   mapp<=25;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=24515;
 end   
19'd66003: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=97;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd66004: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=24;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd66005: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=11;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd66006: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=67;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd66007: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=65;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd66008: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=40;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd66009: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=79;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd66010: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd66011: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=48;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=35541;
 end   
19'd66012: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=4;
   mapp<=28;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=39080;
 end   
19'd66013: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=48;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd66014: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=65;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd66015: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=21;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd66016: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=33;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd66017: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=75;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd66018: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=41;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd66019: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=14;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd66020: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd66021: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd66163: begin  
rid<=1;
end
19'd66164: begin  
end
19'd66165: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd66166: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd66167: begin  
rid<=0;
end
19'd66301: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=21;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16098;
 end   
19'd66302: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=84;
   mapp<=76;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15726;
 end   
19'd66303: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=88;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd66304: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=66;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd66305: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd66306: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=29;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=26237;
 end   
19'd66307: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=89;
   mapp<=80;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=24303;
 end   
19'd66308: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=43;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd66309: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=4;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd66310: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=1;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd66311: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd66453: begin  
rid<=1;
end
19'd66454: begin  
end
19'd66455: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd66456: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd66457: begin  
rid<=0;
end
19'd66601: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=28;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16182;
 end   
19'd66602: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=66;
   mapp<=36;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=17936;
 end   
19'd66603: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=72;
   mapp<=52;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=19126;
 end   
19'd66604: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=93;
   mapp<=82;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=21123;
 end   
19'd66605: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=58;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd66606: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=79;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd66607: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=83;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd66608: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=94;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=31444;
 end   
19'd66609: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=1;
   mapp<=23;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=21470;
 end   
19'd66610: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=53;
   mapp<=97;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=31400;
 end   
19'd66611: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=20;
   mapp<=96;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=31836;
 end   
19'd66612: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=3;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd66613: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=72;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd66614: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=20;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd66615: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd66757: begin  
rid<=1;
end
19'd66758: begin  
end
19'd66759: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd66760: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd66761: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd66762: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd66763: begin  
rid<=0;
end
19'd66901: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=90;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7706;
 end   
19'd66902: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=68;
   mapp<=33;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9442;
 end   
19'd66903: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=26;
   mapp<=57;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12642;
 end   
19'd66904: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=28;
   mapp<=65;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=12012;
 end   
19'd66905: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=32;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=11950;
 end   
19'd66906: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd66907: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd66908: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd66909: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=27;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14378;
 end   
19'd66910: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=10;
   mapp<=44;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=14689;
 end   
19'd66911: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=27;
   mapp<=3;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=14350;
 end   
19'd66912: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=82;
   mapp<=49;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=14566;
 end   
19'd66913: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=33;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=16421;
 end   
19'd66914: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd66915: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd66916: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd66917: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd67059: begin  
rid<=1;
end
19'd67060: begin  
end
19'd67061: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd67062: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd67063: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd67064: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd67065: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd67066: begin  
rid<=0;
end
19'd67201: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=18;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13100;
 end   
19'd67202: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=81;
   mapp<=61;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=16526;
 end   
19'd67203: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=58;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd67204: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=3;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd67205: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=58;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd67206: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd67207: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=22;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=28597;
 end   
19'd67208: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=56;
   mapp<=64;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=36561;
 end   
19'd67209: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=67;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd67210: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=60;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd67211: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=98;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd67212: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=43;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd67213: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd67355: begin  
rid<=1;
end
19'd67356: begin  
end
19'd67357: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd67358: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd67359: begin  
rid<=0;
end
19'd67501: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=98;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5554;
 end   
19'd67502: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=71;
   mapp<=52;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9508;
 end   
19'd67503: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=62;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6877;
 end   
19'd67504: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=11;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1889;
 end   
19'd67505: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=11;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=7721;
 end   
19'd67506: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=93;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=9519;
 end   
19'd67507: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=5;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=6301;
 end   
19'd67508: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=81;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=11629;
 end   
19'd67509: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=51;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=9338;
 end   
19'd67510: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd67511: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=39;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8132;
 end   
19'd67512: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=10;
   mapp<=94;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=14014;
 end   
19'd67513: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=84;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=10503;
 end   
19'd67514: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=35;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=3254;
 end   
19'd67515: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=8271;
 end   
19'd67516: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=55;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=12214;
 end   
19'd67517: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=55;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=8676;
 end   
19'd67518: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=23;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=13026;
 end   
19'd67519: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=50;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=12168;
 end   
19'd67520: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd67521: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd67663: begin  
rid<=1;
end
19'd67664: begin  
end
19'd67665: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd67666: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd67667: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd67668: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd67669: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd67670: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd67671: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd67672: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd67673: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd67674: begin  
rid<=0;
end
19'd67801: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=19;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9847;
 end   
19'd67802: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=48;
   mapp<=10;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9949;
 end   
19'd67803: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=89;
   mapp<=95;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9847;
 end   
19'd67804: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=71;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=12973;
 end   
19'd67805: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=51;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd67806: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=95;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd67807: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=11772;
 end   
19'd67808: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=7;
   mapp<=37;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=15484;
 end   
19'd67809: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=34;
   mapp<=49;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=17510;
 end   
19'd67810: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=84;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=18342;
 end   
19'd67811: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=77;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd67812: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd67813: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd67955: begin  
rid<=1;
end
19'd67956: begin  
end
19'd67957: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd67958: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd67959: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd67960: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd67961: begin  
rid<=0;
end
19'd68101: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=65;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16483;
 end   
19'd68102: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=38;
   mapp<=62;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12177;
 end   
19'd68103: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=45;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd68104: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=28;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd68105: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=94;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd68106: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd68107: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=57;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=21853;
 end   
19'd68108: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=12;
   mapp<=78;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=19009;
 end   
19'd68109: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=1;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd68110: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=99;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd68111: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=27;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd68112: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd68113: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd68255: begin  
rid<=1;
end
19'd68256: begin  
end
19'd68257: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd68258: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd68259: begin  
rid<=0;
end
19'd68401: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=42;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3990;
 end   
19'd68402: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=67;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6375;
 end   
19'd68403: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=76;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7714;
 end   
19'd68404: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=55;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=9070;
 end   
19'd68405: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd68547: begin  
rid<=1;
end
19'd68548: begin  
end
19'd68549: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd68550: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd68551: begin  
rid<=0;
end
19'd68701: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=47;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1236;
 end   
19'd68702: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=73;
   mapp<=15;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1204;
 end   
19'd68703: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=65;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=950;
 end   
19'd68704: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=49;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=732;
 end   
19'd68705: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=37;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1186;
 end   
19'd68706: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=69;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=722;
 end   
19'd68707: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=31;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd68708: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=68;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8752;
 end   
19'd68709: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=52;
   mapp<=53;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8978;
 end   
19'd68710: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=78;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=9378;
 end   
19'd68711: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=56;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=8945;
 end   
19'd68712: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=81;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=11891;
 end   
19'd68713: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=95;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=11930;
 end   
19'd68714: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=86;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd68715: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd68857: begin  
rid<=1;
end
19'd68858: begin  
end
19'd68859: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd68860: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd68861: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd68862: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd68863: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd68864: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd68865: begin  
rid<=0;
end
19'd69001: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=58;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=15982;
 end   
19'd69002: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=38;
   mapp<=59;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10616;
 end   
19'd69003: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=54;
   mapp<=52;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=13880;
 end   
19'd69004: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=72;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd69005: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=8;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd69006: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=56;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd69007: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=74;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=22205;
 end   
19'd69008: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=19;
   mapp<=47;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=13398;
 end   
19'd69009: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=7;
   mapp<=3;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15877;
 end   
19'd69010: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=5;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd69011: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=99;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd69012: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd69013: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd69155: begin  
rid<=1;
end
19'd69156: begin  
end
19'd69157: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd69158: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd69159: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd69160: begin  
rid<=0;
end
19'd69301: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=99;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12514;
 end   
19'd69302: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=54;
   mapp<=92;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=18727;
 end   
19'd69303: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=67;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd69304: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=12;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd69305: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=14;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd69306: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=29;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd69307: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd69308: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=47;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=32386;
 end   
19'd69309: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=99;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=34570;
 end   
19'd69310: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=89;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd69311: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=74;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd69312: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=36;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd69313: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=12;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd69314: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd69315: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd69457: begin  
rid<=1;
end
19'd69458: begin  
end
19'd69459: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd69460: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd69461: begin  
rid<=0;
end
19'd69601: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=91;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=273;
 end   
19'd69602: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=29;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=2651;
 end   
19'd69603: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd69745: begin  
rid<=1;
end
19'd69746: begin  
end
19'd69747: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd69748: begin  
rid<=0;
end
19'd69901: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=96;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4992;
 end   
19'd69902: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=46;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2402;
 end   
19'd69903: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=83;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4336;
 end   
19'd69904: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=97;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5074;
 end   
19'd69905: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=54;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2848;
 end   
19'd69906: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=32;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=1714;
 end   
19'd69907: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=2;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=164;
 end   
19'd69908: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=45;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=2410;
 end   
19'd69909: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=24;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=6816;
 end   
19'd69910: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=81;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8558;
 end   
19'd69911: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=95;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=11556;
 end   
19'd69912: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=23;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6822;
 end   
19'd69913: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=32;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=5280;
 end   
19'd69914: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=43;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=4982;
 end   
19'd69915: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=2;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=316;
 end   
19'd69916: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=69;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=7654;
 end   
19'd69917: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd70059: begin  
rid<=1;
end
19'd70060: begin  
end
19'd70061: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd70062: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd70063: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd70064: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd70065: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd70066: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd70067: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd70068: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd70069: begin  
rid<=0;
end
19'd70201: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=52;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13475;
 end   
19'd70202: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=99;
   mapp<=99;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12573;
 end   
19'd70203: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=50;
   mapp<=35;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12361;
 end   
19'd70204: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd70205: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd70206: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=90;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=23696;
 end   
19'd70207: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=4;
   mapp<=45;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=22462;
 end   
19'd70208: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=77;
   mapp<=93;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=24788;
 end   
19'd70209: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd70210: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd70211: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd70353: begin  
rid<=1;
end
19'd70354: begin  
end
19'd70355: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd70356: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd70357: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd70358: begin  
rid<=0;
end
19'd70501: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=37;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=20291;
 end   
19'd70502: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=15;
   mapp<=28;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=23788;
 end   
19'd70503: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=89;
   mapp<=28;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=27305;
 end   
19'd70504: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=81;
   mapp<=22;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=28848;
 end   
19'd70505: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=74;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd70506: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=59;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd70507: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=50;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd70508: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd70509: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd70510: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd70511: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=61;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=34797;
 end   
19'd70512: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=46;
   mapp<=60;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=37811;
 end   
19'd70513: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=58;
   mapp<=27;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=40870;
 end   
19'd70514: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=94;
   mapp<=33;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=42699;
 end   
19'd70515: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=71;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd70516: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=45;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd70517: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=2;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd70518: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd70519: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd70520: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd70521: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd70663: begin  
rid<=1;
end
19'd70664: begin  
end
19'd70665: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd70666: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd70667: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd70668: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd70669: begin  
rid<=0;
end
19'd70801: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=35;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14766;
 end   
19'd70802: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=92;
   mapp<=53;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12618;
 end   
19'd70803: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=18;
   mapp<=60;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=13769;
 end   
19'd70804: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=65;
   mapp<=86;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7368;
 end   
19'd70805: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=70;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd70806: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd70807: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd70808: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd70809: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=26;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=20309;
 end   
19'd70810: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=1;
   mapp<=25;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=23158;
 end   
19'd70811: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=73;
   mapp<=46;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=17577;
 end   
19'd70812: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=6;
   mapp<=44;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=15000;
 end   
19'd70813: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=80;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd70814: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd70815: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd70816: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd70817: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd70959: begin  
rid<=1;
end
19'd70960: begin  
end
19'd70961: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd70962: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd70963: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd70964: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd70965: begin  
rid<=0;
end
19'd71101: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=23;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2891;
 end   
19'd71102: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=57;
   mapp<=14;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5197;
 end   
19'd71103: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=706;
 end   
19'd71104: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=49;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4797;
 end   
19'd71105: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=22;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3232;
 end   
19'd71106: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=85;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=8653;
 end   
19'd71107: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=62;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=5730;
 end   
19'd71108: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=2;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=1204;
 end   
19'd71109: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=68;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=7304;
 end   
19'd71110: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=74;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=7552;
 end   
19'd71111: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=52;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd71112: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=38;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=6885;
 end   
19'd71113: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=62;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=9468;
 end   
19'd71114: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=37;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=5002;
 end   
19'd71115: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=72;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=11473;
 end   
19'd71116: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=92;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=7648;
 end   
19'd71117: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=10158;
 end   
19'd71118: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=43;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=8459;
 end   
19'd71119: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=19;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=4951;
 end   
19'd71120: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=81;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=13642;
 end   
19'd71121: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=70;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=14097;
 end   
19'd71122: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=91;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd71123: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd71265: begin  
rid<=1;
end
19'd71266: begin  
end
19'd71267: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd71268: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd71269: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd71270: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd71271: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd71272: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd71273: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd71274: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd71275: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd71276: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd71277: begin  
rid<=0;
end
19'd71401: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=50;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=27009;
 end   
19'd71402: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=93;
   mapp<=85;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=26798;
 end   
19'd71403: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=85;
   mapp<=79;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=24006;
 end   
19'd71404: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=16;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd71405: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=8;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd71406: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=88;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd71407: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=99;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd71408: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=25;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd71409: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=96;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd71410: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=77;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=43111;
 end   
19'd71411: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=98;
   mapp<=31;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=44412;
 end   
19'd71412: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=51;
   mapp<=14;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=39674;
 end   
19'd71413: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=88;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd71414: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=63;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd71415: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=53;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd71416: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=5;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd71417: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=41;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd71418: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=67;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd71419: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd71561: begin  
rid<=1;
end
19'd71562: begin  
end
19'd71563: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd71564: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd71565: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd71566: begin  
rid<=0;
end
19'd71701: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=38;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16131;
 end   
19'd71702: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=21;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=16866;
 end   
19'd71703: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=45;
   mapp<=18;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=15446;
 end   
19'd71704: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=23;
   mapp<=72;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=14324;
 end   
19'd71705: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=43;
   mapp<=94;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=22950;
 end   
19'd71706: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=65;
   mapp<=70;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=26555;
 end   
19'd71707: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=18;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd71708: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=35;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd71709: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd71710: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=99;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd71711: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=99;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd71712: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=22;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=30298;
 end   
19'd71713: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=56;
   mapp<=54;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=30071;
 end   
19'd71714: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=18;
   mapp<=24;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=28624;
 end   
19'd71715: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=75;
   mapp<=31;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=31247;
 end   
19'd71716: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=92;
   mapp<=66;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=36896;
 end   
19'd71717: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=10;
   mapp<=29;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=35278;
 end   
19'd71718: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=61;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd71719: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=32;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd71720: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=28;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd71721: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=22;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd71722: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=49;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd71723: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd71865: begin  
rid<=1;
end
19'd71866: begin  
end
19'd71867: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd71868: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd71869: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd71870: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd71871: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd71872: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd71873: begin  
rid<=0;
end
19'd72001: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=40;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13200;
 end   
19'd72002: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=40;
   mapp<=78;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=14793;
 end   
19'd72003: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=66;
   mapp<=77;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=13134;
 end   
19'd72004: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=81;
   mapp<=38;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=9479;
 end   
19'd72005: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=75;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=9609;
 end   
19'd72006: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=44;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7085;
 end   
19'd72007: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd72008: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd72009: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd72010: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=3;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=19117;
 end   
19'd72011: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=76;
   mapp<=47;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20263;
 end   
19'd72012: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=40;
   mapp<=51;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=16089;
 end   
19'd72013: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=23;
   mapp<=7;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=15087;
 end   
19'd72014: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=51;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=14573;
 end   
19'd72015: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=10;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=14734;
 end   
19'd72016: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd72017: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd72018: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd72019: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd72161: begin  
rid<=1;
end
19'd72162: begin  
end
19'd72163: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd72164: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd72165: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd72166: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd72167: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd72168: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd72169: begin  
rid<=0;
end
19'd72301: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=99;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9669;
 end   
19'd72302: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=48;
   mapp<=6;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9707;
 end   
19'd72303: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=30;
   mapp<=85;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7458;
 end   
19'd72304: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=73;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6775;
 end   
19'd72305: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=58;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=11278;
 end   
19'd72306: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=16;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7863;
 end   
19'd72307: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=84;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=8929;
 end   
19'd72308: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=73;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=5633;
 end   
19'd72309: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=31;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=9298;
 end   
19'd72310: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=4;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd72311: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=83;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd72312: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=87;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=19674;
 end   
19'd72313: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=64;
   mapp<=22;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=17967;
 end   
19'd72314: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=68;
   mapp<=10;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=16504;
 end   
19'd72315: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=94;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=17297;
 end   
19'd72316: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=79;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=19063;
 end   
19'd72317: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=23;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=10724;
 end   
19'd72318: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=9;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=11412;
 end   
19'd72319: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=57;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=12572;
 end   
19'd72320: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=41;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=15669;
 end   
19'd72321: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=85;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd72322: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=77;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd72323: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd72465: begin  
rid<=1;
end
19'd72466: begin  
end
19'd72467: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd72468: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd72469: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd72470: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd72471: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd72472: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd72473: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd72474: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd72475: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd72476: begin  
rid<=0;
end
19'd72601: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=69;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4750;
 end   
19'd72602: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=38;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5039;
 end   
19'd72603: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=4;
   mapp<=49;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7351;
 end   
19'd72604: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=76;
   mapp<=17;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6809;
 end   
19'd72605: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=9;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=7503;
 end   
19'd72606: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=43;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=12663;
 end   
19'd72607: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=67;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=14429;
 end   
19'd72608: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd72609: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd72610: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd72611: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=42;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=18017;
 end   
19'd72612: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=40;
   mapp<=91;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=15262;
 end   
19'd72613: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=89;
   mapp<=93;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=22515;
 end   
19'd72614: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=94;
   mapp<=9;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=22448;
 end   
19'd72615: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=20;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=20373;
 end   
19'd72616: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=97;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=21709;
 end   
19'd72617: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=62;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=23699;
 end   
19'd72618: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd72619: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd72620: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd72621: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd72763: begin  
rid<=1;
end
19'd72764: begin  
end
19'd72765: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd72766: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd72767: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd72768: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd72769: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd72770: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd72771: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd72772: begin  
rid<=0;
end
19'd72901: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=43;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=21588;
 end   
19'd72902: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=66;
   mapp<=46;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=23017;
 end   
19'd72903: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=74;
   mapp<=64;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=20217;
 end   
19'd72904: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=45;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd72905: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=88;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd72906: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=49;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd72907: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=27;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd72908: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=85;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=35917;
 end   
19'd72909: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=14;
   mapp<=4;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=32374;
 end   
19'd72910: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=50;
   mapp<=81;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=31620;
 end   
19'd72911: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=32;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd72912: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=73;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd72913: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=43;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd72914: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd72915: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd73057: begin  
rid<=1;
end
19'd73058: begin  
end
19'd73059: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd73060: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd73061: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd73062: begin  
rid<=0;
end
19'd73201: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=35;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1365;
 end   
19'd73202: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2390;
 end   
19'd73203: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=89;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3135;
 end   
19'd73204: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=83;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=2935;
 end   
19'd73205: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=9;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=355;
 end   
19'd73206: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=87;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=3095;
 end   
19'd73207: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=95;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=3385;
 end   
19'd73208: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=45;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=1645;
 end   
19'd73209: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=12;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=500;
 end   
19'd73210: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=39;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=1455;
 end   
19'd73211: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=77;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5061;
 end   
19'd73212: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=79;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8473;
 end   
19'd73213: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=7;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=3674;
 end   
19'd73214: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=30;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=5245;
 end   
19'd73215: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=54;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=4513;
 end   
19'd73216: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=1;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=3172;
 end   
19'd73217: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=40;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=6465;
 end   
19'd73218: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=43;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=4956;
 end   
19'd73219: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=18;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=1886;
 end   
19'd73220: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=12;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=2379;
 end   
19'd73221: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd73363: begin  
rid<=1;
end
19'd73364: begin  
end
19'd73365: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd73366: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd73367: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd73368: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd73369: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd73370: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd73371: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd73372: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd73373: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd73374: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd73375: begin  
rid<=0;
end
19'd73501: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=57;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8375;
 end   
19'd73502: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=2;
   mapp<=85;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5527;
 end   
19'd73503: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=39;
   mapp<=86;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10783;
 end   
19'd73504: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=6;
   mapp<=20;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=10092;
 end   
19'd73505: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=76;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=13600;
 end   
19'd73506: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=24;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=10344;
 end   
19'd73507: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=52;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=12511;
 end   
19'd73508: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=37;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=14950;
 end   
19'd73509: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=35;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd73510: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=99;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd73511: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd73512: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=75;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=18382;
 end   
19'd73513: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=20;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=14868;
 end   
19'd73514: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=92;
   mapp<=6;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=24918;
 end   
19'd73515: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=65;
   mapp<=21;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=21203;
 end   
19'd73516: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=47;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=22871;
 end   
19'd73517: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=58;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=21987;
 end   
19'd73518: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=84;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=24044;
 end   
19'd73519: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=31;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=20280;
 end   
19'd73520: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=29;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd73521: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=82;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd73522: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=5;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd73523: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd73665: begin  
rid<=1;
end
19'd73666: begin  
end
19'd73667: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd73668: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd73669: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd73670: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd73671: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd73672: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd73673: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd73674: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd73675: begin  
rid<=0;
end
19'd73801: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=80;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10924;
 end   
19'd73802: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=69;
   mapp<=70;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15852;
 end   
19'd73803: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=72;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd73804: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=15;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd73805: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=0;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd73806: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=54;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=23006;
 end   
19'd73807: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=29;
   mapp<=36;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=29386;
 end   
19'd73808: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=82;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd73809: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=51;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd73810: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=0;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd73811: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd73953: begin  
rid<=1;
end
19'd73954: begin  
end
19'd73955: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd73956: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd73957: begin  
rid<=0;
end
19'd74101: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=73;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5097;
 end   
19'd74102: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=61;
   mapp<=76;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7823;
 end   
19'd74103: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=97;
   mapp<=4;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7437;
 end   
19'd74104: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=95;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=2365;
 end   
19'd74105: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=25;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6773;
 end   
19'd74106: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=85;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd74107: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd74108: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=73;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12116;
 end   
19'd74109: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=79;
   mapp<=60;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=11770;
 end   
19'd74110: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=9;
   mapp<=18;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=11850;
 end   
19'd74111: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=62;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6935;
 end   
19'd74112: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=24;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=13385;
 end   
19'd74113: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=74;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd74114: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=82;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd74115: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd74257: begin  
rid<=1;
end
19'd74258: begin  
end
19'd74259: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd74260: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd74261: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd74262: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd74263: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd74264: begin  
rid<=0;
end
19'd74401: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=86;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=22167;
 end   
19'd74402: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=66;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd74403: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=89;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd74404: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=51;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd74405: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=4;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd74406: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=33;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd74407: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=94;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd74408: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=64;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=44309;
 end   
19'd74409: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=16;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd74410: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=14;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd74411: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=66;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd74412: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=96;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd74413: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=73;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd74414: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=48;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd74415: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd74557: begin  
rid<=1;
end
19'd74558: begin  
end
19'd74559: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd74560: begin  
rid<=0;
end
19'd74701: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=89;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5469;
 end   
19'd74702: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=20;
   mapp<=91;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9429;
 end   
19'd74703: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd74704: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=81;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=13332;
 end   
19'd74705: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=71;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=16938;
 end   
19'd74706: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd74707: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd74849: begin  
rid<=1;
end
19'd74850: begin  
end
19'd74851: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd74852: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd74853: begin  
rid<=0;
end
19'd75001: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=30;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5061;
 end   
19'd75002: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=38;
   mapp<=54;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8049;
 end   
19'd75003: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=91;
   mapp<=9;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9246;
 end   
19'd75004: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=39;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6171;
 end   
19'd75005: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=53;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=7104;
 end   
19'd75006: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=48;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7658;
 end   
19'd75007: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=67;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=8560;
 end   
19'd75008: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=54;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=8980;
 end   
19'd75009: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=77;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=11434;
 end   
19'd75010: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=90;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd75011: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=97;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd75012: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=62;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=13742;
 end   
19'd75013: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=36;
   mapp<=73;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20014;
 end   
19'd75014: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=29;
   mapp<=89;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=20765;
 end   
19'd75015: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=88;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=21511;
 end   
19'd75016: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=39;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=19142;
 end   
19'd75017: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=85;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=21374;
 end   
19'd75018: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=41;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=17527;
 end   
19'd75019: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=67;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=19532;
 end   
19'd75020: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=20;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=21117;
 end   
19'd75021: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=60;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd75022: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=47;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd75023: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd75165: begin  
rid<=1;
end
19'd75166: begin  
end
19'd75167: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd75168: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd75169: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd75170: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd75171: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd75172: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd75173: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd75174: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd75175: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd75176: begin  
rid<=0;
end
19'd75301: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=92;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=552;
 end   
19'd75302: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=89;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8198;
 end   
19'd75303: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=84;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7748;
 end   
19'd75304: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=3;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=306;
 end   
19'd75305: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=60;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5560;
 end   
19'd75306: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=62;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=5754;
 end   
19'd75307: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=32;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=3004;
 end   
19'd75308: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=70;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=3562;
 end   
19'd75309: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=63;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12608;
 end   
19'd75310: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=23;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=9358;
 end   
19'd75311: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=11;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=1076;
 end   
19'd75312: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=40;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=8360;
 end   
19'd75313: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=92;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=12194;
 end   
19'd75314: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=43;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=6014;
 end   
19'd75315: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd75457: begin  
rid<=1;
end
19'd75458: begin  
end
19'd75459: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd75460: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd75461: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd75462: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd75463: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd75464: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd75465: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd75466: begin  
rid<=0;
end
19'd75601: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=56;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12208;
 end   
19'd75602: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=3;
   mapp<=76;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10008;
 end   
19'd75603: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=64;
   mapp<=45;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=15304;
 end   
19'd75604: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=98;
   mapp<=86;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=8592;
 end   
19'd75605: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=8;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=9752;
 end   
19'd75606: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=78;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd75607: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd75608: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd75609: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=43;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=15552;
 end   
19'd75610: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=27;
   mapp<=11;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18939;
 end   
19'd75611: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=14;
   mapp<=93;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=17869;
 end   
19'd75612: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=90;
   mapp<=17;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=9974;
 end   
19'd75613: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=16;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=14218;
 end   
19'd75614: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=1;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd75615: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=39;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd75616: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=44;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd75617: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd75759: begin  
rid<=1;
end
19'd75760: begin  
end
19'd75761: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd75762: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd75763: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd75764: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd75765: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd75766: begin  
rid<=0;
end
19'd75901: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=37;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7011;
 end   
19'd75902: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=34;
   mapp<=33;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8561;
 end   
19'd75903: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=77;
   mapp<=40;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10410;
 end   
19'd75904: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=71;
   mapp<=1;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7572;
 end   
19'd75905: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=83;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=8800;
 end   
19'd75906: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd75907: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd75908: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd75909: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=90;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16954;
 end   
19'd75910: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=27;
   mapp<=63;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=22972;
 end   
19'd75911: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=58;
   mapp<=59;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=26566;
 end   
19'd75912: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=71;
   mapp<=40;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=21172;
 end   
19'd75913: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=68;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=24604;
 end   
19'd75914: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd75915: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd75916: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd75917: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd76059: begin  
rid<=1;
end
19'd76060: begin  
end
19'd76061: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd76062: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd76063: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd76064: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd76065: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd76066: begin  
rid<=0;
end
19'd76201: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=88;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7374;
 end   
19'd76202: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=64;
   mapp<=34;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11497;
 end   
19'd76203: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=73;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10211;
 end   
19'd76204: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=55;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=12545;
 end   
19'd76205: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=7;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=9182;
 end   
19'd76206: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=99;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=16157;
 end   
19'd76207: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=30;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=7719;
 end   
19'd76208: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=75;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=9709;
 end   
19'd76209: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=3;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=9702;
 end   
19'd76210: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd76211: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd76212: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=4;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12414;
 end   
19'd76213: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=16;
   mapp<=58;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=17272;
 end   
19'd76214: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=49;
   mapp<=80;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15059;
 end   
19'd76215: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=87;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=14554;
 end   
19'd76216: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=64;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=10283;
 end   
19'd76217: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=13;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=18965;
 end   
19'd76218: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=13;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=12033;
 end   
19'd76219: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=52;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=14859;
 end   
19'd76220: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=70;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=14464;
 end   
19'd76221: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd76222: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd76223: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd76365: begin  
rid<=1;
end
19'd76366: begin  
end
19'd76367: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd76368: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd76369: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd76370: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd76371: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd76372: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd76373: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd76374: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd76375: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd76376: begin  
rid<=0;
end
19'd76501: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=26;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3145;
 end   
19'd76502: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=37;
   mapp<=59;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2728;
 end   
19'd76503: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=32;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2887;
 end   
19'd76504: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=55;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1645;
 end   
19'd76505: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd76506: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=82;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=9047;
 end   
19'd76507: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=35;
   mapp<=14;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=5801;
 end   
19'd76508: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=55;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=10547;
 end   
19'd76509: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=90;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=10635;
 end   
19'd76510: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd76511: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd76653: begin  
rid<=1;
end
19'd76654: begin  
end
19'd76655: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd76656: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd76657: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd76658: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd76659: begin  
rid<=0;
end
19'd76801: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=74;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=20006;
 end   
19'd76802: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=24;
   mapp<=38;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=19697;
 end   
19'd76803: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=44;
   mapp<=56;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=14711;
 end   
19'd76804: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=63;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd76805: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=49;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd76806: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=76;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd76807: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=97;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd76808: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=34;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd76809: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=47;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd76810: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=26;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd76811: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=81;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=41564;
 end   
19'd76812: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=71;
   mapp<=44;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=42475;
 end   
19'd76813: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=68;
   mapp<=92;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=36372;
 end   
19'd76814: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=13;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd76815: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=66;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd76816: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=30;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd76817: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=6;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd76818: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=9;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd76819: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=90;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd76820: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=59;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd76821: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd76963: begin  
rid<=1;
end
19'd76964: begin  
end
19'd76965: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd76966: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd76967: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd76968: begin  
rid<=0;
end
19'd77101: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=96;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11400;
 end   
19'd77102: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=83;
   mapp<=3;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10647;
 end   
19'd77103: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=50;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd77104: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=57;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd77105: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=0;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd77106: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=3;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=19582;
 end   
19'd77107: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=73;
   mapp<=12;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=22893;
 end   
19'd77108: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=91;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd77109: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=16;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd77110: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=0;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd77111: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd77253: begin  
rid<=1;
end
19'd77254: begin  
end
19'd77255: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd77256: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd77257: begin  
rid<=0;
end
19'd77401: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=43;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=774;
 end   
19'd77402: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=88;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1594;
 end   
19'd77403: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=97;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1766;
 end   
19'd77404: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=11;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=228;
 end   
19'd77405: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=91;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1678;
 end   
19'd77406: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=74;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=1382;
 end   
19'd77407: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=25;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=2349;
 end   
19'd77408: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=7;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=2035;
 end   
19'd77409: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=70;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=6176;
 end   
19'd77410: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=21;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=1551;
 end   
19'd77411: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=27;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=3379;
 end   
19'd77412: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=58;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=5036;
 end   
19'd77413: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd77555: begin  
rid<=1;
end
19'd77556: begin  
end
19'd77557: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd77558: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd77559: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd77560: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd77561: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd77562: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd77563: begin  
rid<=0;
end
19'd77701: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=11;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5282;
 end   
19'd77702: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=12;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd77703: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=9;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd77704: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=35;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd77705: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=63;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd77706: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=88;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=15738;
 end   
19'd77707: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=39;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd77708: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=5;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd77709: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=70;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd77710: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=40;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd77711: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd77853: begin  
rid<=1;
end
19'd77854: begin  
end
19'd77855: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd77856: begin  
rid<=0;
end
19'd78001: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=37;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1036;
 end   
19'd78002: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=0;
   mapp<=85;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3155;
 end   
19'd78003: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=97;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=2976;
 end   
19'd78004: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=0;
   mapp<=24;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=5483;
 end   
19'd78005: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd78147: begin  
rid<=1;
end
19'd78148: begin  
end
19'd78149: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd78150: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd78151: begin  
rid<=0;
end
19'd78301: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=2;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8017;
 end   
19'd78302: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=14;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd78303: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=29;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd78304: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=94;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd78305: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=26;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd78306: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=99;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=23490;
 end   
19'd78307: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=3;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd78308: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=42;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd78309: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=80;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd78310: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=16;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd78311: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd78453: begin  
rid<=1;
end
19'd78454: begin  
end
19'd78455: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd78456: begin  
rid<=0;
end
19'd78601: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=30;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1740;
 end   
19'd78602: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=53;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3084;
 end   
19'd78603: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=51;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2978;
 end   
19'd78604: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=62;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3626;
 end   
19'd78605: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=44;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2592;
 end   
19'd78606: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=49;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=2892;
 end   
19'd78607: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=85;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=4990;
 end   
19'd78608: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=72;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5700;
 end   
19'd78609: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=89;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=7979;
 end   
19'd78610: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=58;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=6168;
 end   
19'd78611: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=52;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6486;
 end   
19'd78612: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=29;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=4187;
 end   
19'd78613: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=40;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=5092;
 end   
19'd78614: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=60;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=8290;
 end   
19'd78615: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd78757: begin  
rid<=1;
end
19'd78758: begin  
end
19'd78759: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd78760: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd78761: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd78762: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd78763: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd78764: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd78765: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd78766: begin  
rid<=0;
end
19'd78901: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=56;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11744;
 end   
19'd78902: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=51;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd78903: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=91;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd78904: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=34;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd78905: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=31;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd78906: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=22;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd78907: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=29;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=23532;
 end   
19'd78908: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=85;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd78909: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=2;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd78910: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=10;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd78911: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=27;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd78912: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=74;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd78913: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd79055: begin  
rid<=1;
end
19'd79056: begin  
end
19'd79057: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd79058: begin  
rid<=0;
end
19'd79201: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=98;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4116;
 end   
19'd79202: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=55;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5400;
 end   
19'd79203: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=93;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9134;
 end   
19'd79204: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=65;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6400;
 end   
19'd79205: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=28;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2784;
 end   
19'd79206: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=72;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7106;
 end   
19'd79207: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=84;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=8292;
 end   
19'd79208: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=26;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=2618;
 end   
19'd79209: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=78;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5910;
 end   
19'd79210: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=1;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=5478;
 end   
19'd79211: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=87;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15920;
 end   
19'd79212: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=88;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=13264;
 end   
19'd79213: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=97;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=10350;
 end   
19'd79214: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=52;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=11162;
 end   
19'd79215: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=75;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=14142;
 end   
19'd79216: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=50;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=6518;
 end   
19'd79217: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd79359: begin  
rid<=1;
end
19'd79360: begin  
end
19'd79361: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd79362: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd79363: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd79364: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd79365: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd79366: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd79367: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd79368: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd79369: begin  
rid<=0;
end
19'd79501: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=21;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7181;
 end   
19'd79502: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=27;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd79503: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=64;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd79504: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=40;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd79505: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=13;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd79506: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=88;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=22124;
 end   
19'd79507: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=21;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd79508: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=64;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd79509: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=3;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd79510: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=54;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd79511: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd79653: begin  
rid<=1;
end
19'd79654: begin  
end
19'd79655: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd79656: begin  
rid<=0;
end
19'd79801: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=2;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6891;
 end   
19'd79802: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=20;
   mapp<=86;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11070;
 end   
19'd79803: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=59;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd79804: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=88;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd79805: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=82;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd79806: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=41;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd79807: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=52;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17011;
 end   
19'd79808: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=50;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18486;
 end   
19'd79809: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=16;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd79810: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=26;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd79811: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=86;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd79812: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=2;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd79813: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd79955: begin  
rid<=1;
end
19'd79956: begin  
end
19'd79957: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd79958: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd79959: begin  
rid<=0;
end
19'd80101: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=81;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8659;
 end   
19'd80102: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=43;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd80103: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=10;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd80104: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=8;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd80105: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=89;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd80106: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=87;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=23539;
 end   
19'd80107: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=71;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd80108: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=90;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd80109: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=72;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd80110: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=18;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd80111: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd80253: begin  
rid<=1;
end
19'd80254: begin  
end
19'd80255: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd80256: begin  
rid<=0;
end
19'd80401: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=4;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8762;
 end   
19'd80402: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=85;
   mapp<=62;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8847;
 end   
19'd80403: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=33;
   mapp<=96;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3192;
 end   
19'd80404: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=13;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4912;
 end   
19'd80405: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd80406: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd80407: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=72;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=15082;
 end   
19'd80408: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=21;
   mapp<=4;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12244;
 end   
19'd80409: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=44;
   mapp<=37;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=10665;
 end   
19'd80410: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=53;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=11944;
 end   
19'd80411: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd80412: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd80413: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd80555: begin  
rid<=1;
end
19'd80556: begin  
end
19'd80557: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd80558: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd80559: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd80560: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd80561: begin  
rid<=0;
end
19'd80701: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=23;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6224;
 end   
19'd80702: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=1;
   mapp<=29;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2494;
 end   
19'd80703: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=43;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd80704: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd80705: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=13;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8855;
 end   
19'd80706: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=53;
   mapp<=31;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=3425;
 end   
19'd80707: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=11;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd80708: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd80709: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd80851: begin  
rid<=1;
end
19'd80852: begin  
end
19'd80853: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd80854: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd80855: begin  
rid<=0;
end
19'd81001: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=16;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4350;
 end   
19'd81002: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=12;
   mapp<=14;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5949;
 end   
19'd81003: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=34;
   mapp<=99;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7588;
 end   
19'd81004: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=49;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4445;
 end   
19'd81005: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=52;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6919;
 end   
19'd81006: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=12;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=2127;
 end   
19'd81007: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=41;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd81008: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=9;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd81009: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=35;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=15545;
 end   
19'd81010: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=62;
   mapp<=80;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=15008;
 end   
19'd81011: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=65;
   mapp<=69;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=12891;
 end   
19'd81012: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=11;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=7114;
 end   
19'd81013: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=17;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=12996;
 end   
19'd81014: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=11;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=9166;
 end   
19'd81015: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=63;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd81016: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=21;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd81017: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd81159: begin  
rid<=1;
end
19'd81160: begin  
end
19'd81161: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd81162: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd81163: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd81164: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd81165: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd81166: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd81167: begin  
rid<=0;
end
19'd81301: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=64;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8944;
 end   
19'd81302: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=42;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd81303: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=44;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd81304: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=25;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=11999;
 end   
19'd81305: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=59;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd81306: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=53;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd81307: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd81449: begin  
rid<=1;
end
19'd81450: begin  
end
19'd81451: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd81452: begin  
rid<=0;
end
19'd81601: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=20;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=23316;
 end   
19'd81602: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=15;
   mapp<=29;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=24658;
 end   
19'd81603: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=44;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd81604: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=78;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd81605: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=58;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd81606: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=84;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd81607: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=38;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd81608: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=83;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd81609: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd81610: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=52;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=33029;
 end   
19'd81611: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=4;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=31928;
 end   
19'd81612: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=46;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd81613: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=12;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd81614: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=4;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd81615: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=45;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd81616: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=25;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd81617: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=44;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd81618: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=49;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd81619: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd81761: begin  
rid<=1;
end
19'd81762: begin  
end
19'd81763: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd81764: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd81765: begin  
rid<=0;
end
19'd81901: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=9;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=288;
 end   
19'd81902: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=16;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=522;
 end   
19'd81903: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=29;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=948;
 end   
19'd81904: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=61;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1982;
 end   
19'd81905: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=33;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1096;
 end   
19'd81906: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=46;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=1668;
 end   
19'd81907: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=32;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=1482;
 end   
19'd81908: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=83;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=3438;
 end   
19'd81909: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=73;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=4172;
 end   
19'd81910: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=39;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=2266;
 end   
19'd81911: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd82053: begin  
rid<=1;
end
19'd82054: begin  
end
19'd82055: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd82056: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd82057: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd82058: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd82059: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd82060: begin  
rid<=0;
end
19'd82201: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=89;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9773;
 end   
19'd82202: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=29;
   mapp<=70;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6733;
 end   
19'd82203: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=60;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd82204: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=89;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17753;
 end   
19'd82205: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=63;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12324;
 end   
19'd82206: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=44;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd82207: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd82349: begin  
rid<=1;
end
19'd82350: begin  
end
19'd82351: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd82352: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd82353: begin  
rid<=0;
end
19'd82501: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=46;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=25317;
 end   
19'd82502: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=43;
   mapp<=13;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=21768;
 end   
19'd82503: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=37;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd82504: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=31;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd82505: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=55;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd82506: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=51;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd82507: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=51;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd82508: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=90;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd82509: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=52;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd82510: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=95;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd82511: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=20;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd82512: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=79;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=48423;
 end   
19'd82513: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=60;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=46921;
 end   
19'd82514: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=15;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd82515: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=9;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd82516: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=72;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd82517: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=61;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd82518: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=52;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd82519: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=70;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd82520: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=23;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd82521: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=64;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd82522: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd82523: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd82665: begin  
rid<=1;
end
19'd82666: begin  
end
19'd82667: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd82668: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd82669: begin  
rid<=0;
end
19'd82801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=83;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16273;
 end   
19'd82802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=33;
   mapp<=78;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15183;
 end   
19'd82803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=95;
   mapp<=43;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=14815;
 end   
19'd82804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=9;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd82805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=72;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd82806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd82807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd82808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=42;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=28768;
 end   
19'd82809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=44;
   mapp<=3;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=26891;
 end   
19'd82810: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=55;
   mapp<=64;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=28256;
 end   
19'd82811: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=59;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd82812: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=68;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd82813: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd82814: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd82815: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd82957: begin  
rid<=1;
end
19'd82958: begin  
end
19'd82959: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd82960: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd82961: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd82962: begin  
rid<=0;
end
19'd83101: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=40;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11060;
 end   
19'd83102: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=25;
   mapp<=47;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10264;
 end   
19'd83103: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=24;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd83104: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=46;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd83105: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd83106: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=38;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd83107: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=31;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd83108: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=21;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd83109: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd83110: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=19;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=31495;
 end   
19'd83111: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=74;
   mapp<=24;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=31918;
 end   
19'd83112: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=87;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd83113: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=30;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd83114: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=45;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd83115: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=16;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd83116: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=44;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd83117: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=99;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd83118: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd83119: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd83261: begin  
rid<=1;
end
19'd83262: begin  
end
19'd83263: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd83264: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd83265: begin  
rid<=0;
end
19'd83401: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=33;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2894;
 end   
19'd83402: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=52;
   mapp<=21;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3126;
 end   
19'd83403: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=11;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd83404: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=29;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd83405: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=24;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd83406: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd83407: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=91;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=24654;
 end   
19'd83408: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=97;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=23355;
 end   
19'd83409: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=13;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd83410: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=71;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd83411: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=86;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd83412: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd83413: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd83555: begin  
rid<=1;
end
19'd83556: begin  
end
19'd83557: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd83558: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd83559: begin  
rid<=0;
end
19'd83701: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=79;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=17583;
 end   
19'd83702: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=98;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd83703: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=67;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd83704: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=45;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd83705: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=3;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd83706: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=30;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd83707: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=20;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd83708: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=25;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd83709: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=34;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd83710: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=21;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd83711: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=33;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd83712: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=86;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=43977;
 end   
19'd83713: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=95;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd83714: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=8;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd83715: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=53;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd83716: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=97;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd83717: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=92;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd83718: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=21;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd83719: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=19;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd83720: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=7;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd83721: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=71;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd83722: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=22;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd83723: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd83865: begin  
rid<=1;
end
19'd83866: begin  
end
19'd83867: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd83868: begin  
rid<=0;
end
19'd84001: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=65;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3380;
 end   
19'd84002: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=51;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3325;
 end   
19'd84003: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=23;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1515;
 end   
19'd84004: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=65;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7020;
 end   
19'd84005: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=80;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8525;
 end   
19'd84006: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=61;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=5480;
 end   
19'd84007: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd84149: begin  
rid<=1;
end
19'd84150: begin  
end
19'd84151: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd84152: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd84153: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd84154: begin  
rid<=0;
end
19'd84301: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=53;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1904;
 end   
19'd84302: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=12;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3216;
 end   
19'd84303: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=82;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd84304: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=89;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=13912;
 end   
19'd84305: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=92;
   mapp<=57;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=15851;
 end   
19'd84306: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=99;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd84307: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd84449: begin  
rid<=1;
end
19'd84450: begin  
end
19'd84451: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd84452: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd84453: begin  
rid<=0;
end
19'd84601: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=20;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10493;
 end   
19'd84602: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=45;
   mapp<=31;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11955;
 end   
19'd84603: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=29;
   mapp<=60;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9738;
 end   
19'd84604: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=68;
   mapp<=0;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=14731;
 end   
19'd84605: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=41;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd84606: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=62;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd84607: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd84608: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=33;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd84609: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd84610: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=36;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=23734;
 end   
19'd84611: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=65;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=25739;
 end   
19'd84612: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=33;
   mapp<=60;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=20549;
 end   
19'd84613: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=29;
   mapp<=64;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=31236;
 end   
19'd84614: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=27;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd84615: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=54;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd84616: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=28;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd84617: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=19;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd84618: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=84;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd84619: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd84761: begin  
rid<=1;
end
19'd84762: begin  
end
19'd84763: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd84764: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd84765: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd84766: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd84767: begin  
rid<=0;
end
19'd84901: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=90;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16884;
 end   
19'd84902: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=69;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd84903: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=44;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd84904: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=99;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd84905: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=43;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd84906: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=55;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd84907: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=64;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd84908: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=29;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=33980;
 end   
19'd84909: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=87;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd84910: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=80;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd84911: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=85;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd84912: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=64;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd84913: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=34;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd84914: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=76;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd84915: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd85057: begin  
rid<=1;
end
19'd85058: begin  
end
19'd85059: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd85060: begin  
rid<=0;
end
19'd85201: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=48;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4032;
 end   
19'd85202: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=0;
   mapp<=47;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2266;
 end   
19'd85203: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=32;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5536;
 end   
19'd85204: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=0;
   mapp<=55;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=4026;
 end   
19'd85205: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd85347: begin  
rid<=1;
end
19'd85348: begin  
end
19'd85349: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd85350: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd85351: begin  
rid<=0;
end
19'd85501: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=4;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10287;
 end   
19'd85502: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=29;
   mapp<=96;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11550;
 end   
19'd85503: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=15;
   mapp<=59;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5932;
 end   
19'd85504: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=65;
   mapp<=24;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5907;
 end   
19'd85505: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=50;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd85506: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd85507: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd85508: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd85509: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=3;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=19892;
 end   
19'd85510: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=6;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20385;
 end   
19'd85511: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=20;
   mapp<=19;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=14667;
 end   
19'd85512: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=70;
   mapp<=96;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=12658;
 end   
19'd85513: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=49;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd85514: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd85515: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd85516: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd85517: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd85659: begin  
rid<=1;
end
19'd85660: begin  
end
19'd85661: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd85662: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd85663: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd85664: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd85665: begin  
rid<=0;
end
19'd85801: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=85;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14949;
 end   
19'd85802: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=63;
   mapp<=87;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15590;
 end   
19'd85803: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=11;
   mapp<=84;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=15884;
 end   
19'd85804: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=66;
   mapp<=29;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=10848;
 end   
19'd85805: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=39;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=12840;
 end   
19'd85806: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=98;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=14387;
 end   
19'd85807: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=73;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=8956;
 end   
19'd85808: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=38;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=6973;
 end   
19'd85809: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd85810: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd85811: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd85812: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=2;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=21067;
 end   
19'd85813: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=48;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20173;
 end   
19'd85814: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=13;
   mapp<=30;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=22262;
 end   
19'd85815: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=26;
   mapp<=65;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=16786;
 end   
19'd85816: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=82;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=18253;
 end   
19'd85817: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=82;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=18834;
 end   
19'd85818: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=31;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=12180;
 end   
19'd85819: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=35;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=12975;
 end   
19'd85820: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd85821: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd85822: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd85823: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd85965: begin  
rid<=1;
end
19'd85966: begin  
end
19'd85967: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd85968: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd85969: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd85970: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd85971: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd85972: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd85973: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd85974: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd85975: begin  
rid<=0;
end
19'd86101: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=70;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11182;
 end   
19'd86102: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=83;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11512;
 end   
19'd86103: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=45;
   mapp<=7;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6871;
 end   
19'd86104: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=28;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd86105: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=59;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd86106: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd86107: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd86108: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=5;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=22341;
 end   
19'd86109: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=47;
   mapp<=21;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20282;
 end   
19'd86110: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=13;
   mapp<=37;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=19463;
 end   
19'd86111: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=86;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd86112: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=84;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd86113: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd86114: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd86115: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd86257: begin  
rid<=1;
end
19'd86258: begin  
end
19'd86259: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd86260: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd86261: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd86262: begin  
rid<=0;
end
19'd86401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=83;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=15348;
 end   
19'd86402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=27;
   mapp<=70;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=21704;
 end   
19'd86403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=99;
   mapp<=39;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=22594;
 end   
19'd86404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=61;
   mapp<=57;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=25606;
 end   
19'd86405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=90;
   mapp<=68;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=23203;
 end   
19'd86406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=56;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=20413;
 end   
19'd86407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=85;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=16940;
 end   
19'd86408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd86409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd86410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd86411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd86412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=99;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=26415;
 end   
19'd86413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=1;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=24479;
 end   
19'd86414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=7;
   mapp<=79;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=39460;
 end   
19'd86415: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=95;
   mapp<=73;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=37880;
 end   
19'd86416: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=19;
   mapp<=6;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=25736;
 end   
19'd86417: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=85;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=33895;
 end   
19'd86418: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=45;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=30092;
 end   
19'd86419: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd86420: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd86421: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd86422: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd86423: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd86565: begin  
rid<=1;
end
19'd86566: begin  
end
19'd86567: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd86568: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd86569: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd86570: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd86571: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd86572: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd86573: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd86574: begin  
rid<=0;
end
19'd86701: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=3;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12579;
 end   
19'd86702: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=88;
   mapp<=60;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=16793;
 end   
19'd86703: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=98;
   mapp<=33;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12395;
 end   
19'd86704: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=75;
   mapp<=52;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=13107;
 end   
19'd86705: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=69;
   mapp<=0;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=9281;
 end   
19'd86706: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=4;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=10053;
 end   
19'd86707: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=90;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd86708: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=43;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd86709: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=57;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd86710: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=57;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd86711: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=98;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=26210;
 end   
19'd86712: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=67;
   mapp<=75;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=32791;
 end   
19'd86713: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=46;
   mapp<=49;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=28700;
 end   
19'd86714: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=9;
   mapp<=90;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=30761;
 end   
19'd86715: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=80;
   mapp<=46;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=22199;
 end   
19'd86716: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=79;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=21430;
 end   
19'd86717: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=81;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd86718: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=7;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd86719: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=19;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd86720: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd86721: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd86863: begin  
rid<=1;
end
19'd86864: begin  
end
19'd86865: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd86866: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd86867: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd86868: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd86869: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd86870: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd86871: begin  
rid<=0;
end
19'd87001: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=64;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11321;
 end   
19'd87002: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=9;
   mapp<=14;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6557;
 end   
19'd87003: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=3;
   mapp<=10;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5831;
 end   
19'd87004: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=44;
   mapp<=55;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7342;
 end   
19'd87005: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=50;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd87006: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=41;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd87007: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd87008: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd87009: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd87010: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=40;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17467;
 end   
19'd87011: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=31;
   mapp<=44;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=15996;
 end   
19'd87012: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=70;
   mapp<=27;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15155;
 end   
19'd87013: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=54;
   mapp<=41;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=20507;
 end   
19'd87014: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=35;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd87015: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=3;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd87016: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd87017: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd87018: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd87019: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd87161: begin  
rid<=1;
end
19'd87162: begin  
end
19'd87163: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd87164: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd87165: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd87166: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd87167: begin  
rid<=0;
end
19'd87301: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=32;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8477;
 end   
19'd87302: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=35;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8048;
 end   
19'd87303: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=17;
   mapp<=17;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12424;
 end   
19'd87304: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=45;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd87305: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=21;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd87306: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=18;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd87307: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=5;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd87308: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=33;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd87309: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=21;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd87310: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=46;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd87311: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd87312: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=42;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=35441;
 end   
19'd87313: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=54;
   mapp<=94;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=29135;
 end   
19'd87314: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=18;
   mapp<=8;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=38861;
 end   
19'd87315: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=90;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd87316: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=24;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd87317: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=79;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd87318: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=65;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd87319: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=54;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd87320: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=71;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd87321: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=22;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd87322: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=44;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd87323: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd87465: begin  
rid<=1;
end
19'd87466: begin  
end
19'd87467: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd87468: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd87469: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd87470: begin  
rid<=0;
end
19'd87601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=41;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9980;
 end   
19'd87602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=17;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=13883;
 end   
19'd87603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=68;
   mapp<=52;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=14951;
 end   
19'd87604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=65;
   mapp<=74;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=15519;
 end   
19'd87605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=77;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=12271;
 end   
19'd87606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=97;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=12360;
 end   
19'd87607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd87608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd87609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd87610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=82;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16601;
 end   
19'd87611: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=35;
   mapp<=55;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=23531;
 end   
19'd87612: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=92;
   mapp<=27;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=26586;
 end   
19'd87613: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=35;
   mapp<=14;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=24096;
 end   
19'd87614: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=83;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=25031;
 end   
19'd87615: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=37;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=23192;
 end   
19'd87616: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd87617: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd87618: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd87619: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd87761: begin  
rid<=1;
end
19'd87762: begin  
end
19'd87763: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd87764: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd87765: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd87766: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd87767: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd87768: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd87769: begin  
rid<=0;
end
19'd87901: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=60;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7978;
 end   
19'd87902: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=65;
   mapp<=28;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11065;
 end   
19'd87903: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=30;
   mapp<=88;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10061;
 end   
19'd87904: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=64;
   mapp<=24;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5437;
 end   
19'd87905: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=23;
   mapp<=34;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6421;
 end   
19'd87906: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=33;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6269;
 end   
19'd87907: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd87908: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd87909: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd87910: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd87911: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=19;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16036;
 end   
19'd87912: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=51;
   mapp<=86;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20070;
 end   
19'd87913: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=41;
   mapp<=8;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=16373;
 end   
19'd87914: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=15;
   mapp<=38;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=15507;
 end   
19'd87915: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=76;
   mapp<=31;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=17109;
 end   
19'd87916: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=65;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=18245;
 end   
19'd87917: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd87918: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd87919: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd87920: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd87921: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd88063: begin  
rid<=1;
end
19'd88064: begin  
end
19'd88065: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd88066: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd88067: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd88068: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd88069: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd88070: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd88071: begin  
rid<=0;
end
19'd88201: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=52;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14797;
 end   
19'd88202: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=30;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd88203: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=74;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd88204: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=81;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd88205: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=42;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd88206: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=80;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=20011;
 end   
19'd88207: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=90;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd88208: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd88209: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=99;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd88210: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=68;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd88211: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd88353: begin  
rid<=1;
end
19'd88354: begin  
end
19'd88355: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd88356: begin  
rid<=0;
end
19'd88501: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=44;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2772;
 end   
19'd88502: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=8;
   mapp<=44;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=450;
 end   
19'd88503: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=856;
 end   
19'd88504: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=19;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1867;
 end   
19'd88505: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=18;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3186;
 end   
19'd88506: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=49;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=4813;
 end   
19'd88507: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=47;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=6165;
 end   
19'd88508: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=80;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=8826;
 end   
19'd88509: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=99;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=7637;
 end   
19'd88510: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=48;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=6426;
 end   
19'd88511: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=84;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd88512: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=40;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=6348;
 end   
19'd88513: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=88;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=4362;
 end   
19'd88514: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=70;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=5290;
 end   
19'd88515: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=97;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=4766;
 end   
19'd88516: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=33;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=5093;
 end   
19'd88517: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=40;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=6277;
 end   
19'd88518: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=22;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=8023;
 end   
19'd88519: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=45;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=10961;
 end   
19'd88520: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=40;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=9261;
 end   
19'd88521: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=27;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=8539;
 end   
19'd88522: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=50;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd88523: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd88665: begin  
rid<=1;
end
19'd88666: begin  
end
19'd88667: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd88668: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd88669: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd88670: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd88671: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd88672: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd88673: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd88674: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd88675: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd88676: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd88677: begin  
rid<=0;
end
19'd88801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=51;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=19602;
 end   
19'd88802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=82;
   mapp<=50;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=20725;
 end   
19'd88803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=39;
   mapp<=30;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=18900;
 end   
19'd88804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=67;
   mapp<=96;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=19138;
 end   
19'd88805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=70;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd88806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=76;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd88807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=43;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd88808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=56;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd88809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=73;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd88810: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd88811: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=98;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=38780;
 end   
19'd88812: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=71;
   mapp<=86;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=39707;
 end   
19'd88813: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=37;
   mapp<=66;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=33725;
 end   
19'd88814: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=61;
   mapp<=33;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=32402;
 end   
19'd88815: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=9;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd88816: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=20;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd88817: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=86;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd88818: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=27;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd88819: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=41;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd88820: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=53;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd88821: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd88963: begin  
rid<=1;
end
19'd88964: begin  
end
19'd88965: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd88966: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd88967: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd88968: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd88969: begin  
rid<=0;
end
19'd89101: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=99;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16866;
 end   
19'd89102: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=81;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd89103: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=71;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=19279;
 end   
19'd89104: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=78;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd89105: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd89247: begin  
rid<=1;
end
19'd89248: begin  
end
19'd89249: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd89250: begin  
rid<=0;
end
19'd89401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=47;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4385;
 end   
19'd89402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=13;
   mapp<=34;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4417;
 end   
19'd89403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=22;
   mapp<=66;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7600;
 end   
19'd89404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=45;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=10739;
 end   
19'd89405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=74;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=8406;
 end   
19'd89406: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=88;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=10544;
 end   
19'd89407: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=22;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=5098;
 end   
19'd89408: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=77;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=10275;
 end   
19'd89409: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=19;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd89410: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=83;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd89411: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=46;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=11395;
 end   
19'd89412: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=24;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=14572;
 end   
19'd89413: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=41;
   mapp<=94;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=19963;
 end   
19'd89414: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=89;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=26221;
 end   
19'd89415: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=98;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=21563;
 end   
19'd89416: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=97;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=22916;
 end   
19'd89417: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=66;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=18308;
 end   
19'd89418: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=60;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=21552;
 end   
19'd89419: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=91;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd89420: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=73;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd89421: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd89563: begin  
rid<=1;
end
19'd89564: begin  
end
19'd89565: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd89566: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd89567: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd89568: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd89569: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd89570: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd89571: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd89572: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd89573: begin  
rid<=0;
end
19'd89701: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=38;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=228;
 end   
19'd89702: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=96;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=586;
 end   
19'd89703: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=18;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=128;
 end   
19'd89704: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=62;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=402;
 end   
19'd89705: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=44;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=304;
 end   
19'd89706: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=26;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=206;
 end   
19'd89707: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=15;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=150;
 end   
19'd89708: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=93;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=628;
 end   
19'd89709: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=69;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=1815;
 end   
19'd89710: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=24;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=1138;
 end   
19'd89711: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=18;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=542;
 end   
19'd89712: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=69;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=1989;
 end   
19'd89713: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=72;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=1960;
 end   
19'd89714: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=70;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=1816;
 end   
19'd89715: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=61;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=1553;
 end   
19'd89716: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=15;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=973;
 end   
19'd89717: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd89859: begin  
rid<=1;
end
19'd89860: begin  
end
19'd89861: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd89862: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd89863: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd89864: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd89865: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd89866: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd89867: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd89868: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd89869: begin  
rid<=0;
end
19'd90001: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=94;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14138;
 end   
19'd90002: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=61;
   mapp<=37;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=13881;
 end   
19'd90003: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=3;
   mapp<=95;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10927;
 end   
19'd90004: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=92;
   mapp<=30;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5931;
 end   
19'd90005: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd90006: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd90007: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd90008: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=61;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=21246;
 end   
19'd90009: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=51;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=22558;
 end   
19'd90010: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=10;
   mapp<=6;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15649;
 end   
19'd90011: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=77;
   mapp<=13;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=14868;
 end   
19'd90012: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd90013: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd90014: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd90015: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd90157: begin  
rid<=1;
end
19'd90158: begin  
end
19'd90159: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd90160: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd90161: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd90162: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd90163: begin  
rid<=0;
end
19'd90301: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=20;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=440;
 end   
19'd90302: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=50;
 end   
19'd90303: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=24;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=500;
 end   
19'd90304: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=96;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1950;
 end   
19'd90305: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=49;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1020;
 end   
19'd90306: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=23;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=510;
 end   
19'd90307: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=12;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=300;
 end   
19'd90308: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=23;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=530;
 end   
19'd90309: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=14;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=360;
 end   
19'd90310: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=71;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=1510;
 end   
19'd90311: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=8;
   pp<=100;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[10]<=260;
 end   
19'd90312: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=4;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=764;
 end   
19'd90313: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=274;
 end   
19'd90314: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=98;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=892;
 end   
19'd90315: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=49;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=2146;
 end   
19'd90316: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=45;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=1200;
 end   
19'd90317: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=97;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=898;
 end   
19'd90318: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=66;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=564;
 end   
19'd90319: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=43;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=702;
 end   
19'd90320: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=48;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=552;
 end   
19'd90321: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=92;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=1878;
 end   
19'd90322: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=31;
   pp<=100;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[10]<=384;
 end   
19'd90323: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd90465: begin  
rid<=1;
end
19'd90466: begin  
end
19'd90467: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd90468: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd90469: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd90470: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd90471: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd90472: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd90473: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd90474: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd90475: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd90476: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd90477: begin  
check0<=expctdoutput[10]-outcheck0;
end
19'd90478: begin  
rid<=0;
end
19'd90601: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=75;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12912;
 end   
19'd90602: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=45;
   mapp<=49;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=16018;
 end   
19'd90603: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=84;
   mapp<=51;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=17207;
 end   
19'd90604: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=33;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd90605: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd90606: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd90607: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=31;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=36457;
 end   
19'd90608: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=99;
   mapp<=99;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=35892;
 end   
19'd90609: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=98;
   mapp<=67;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=32803;
 end   
19'd90610: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=74;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd90611: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd90612: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd90613: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd90755: begin  
rid<=1;
end
19'd90756: begin  
end
19'd90757: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd90758: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd90759: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd90760: begin  
rid<=0;
end
19'd90901: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=45;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2790;
 end   
19'd90902: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=59;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=4501;
 end   
19'd90903: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd91045: begin  
rid<=1;
end
19'd91046: begin  
end
19'd91047: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd91048: begin  
rid<=0;
end
19'd91201: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=96;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=27397;
 end   
19'd91202: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=17;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=20497;
 end   
19'd91203: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=11;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd91204: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=68;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd91205: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=48;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd91206: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=81;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd91207: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=33;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd91208: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=74;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd91209: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd91210: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=11;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=37098;
 end   
19'd91211: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=22;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=31773;
 end   
19'd91212: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=51;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd91213: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd91214: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=42;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd91215: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=30;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd91216: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=25;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd91217: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=30;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd91218: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=51;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd91219: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd91361: begin  
rid<=1;
end
19'd91362: begin  
end
19'd91363: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd91364: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd91365: begin  
rid<=0;
end
19'd91501: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=5;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5415;
 end   
19'd91502: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=66;
   mapp<=80;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=740;
 end   
19'd91503: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=5;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5457;
 end   
19'd91504: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=82;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=2090;
 end   
19'd91505: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=25;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1089;
 end   
19'd91506: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=14;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=912;
 end   
19'd91507: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=12;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=384;
 end   
19'd91508: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=4;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=6162;
 end   
19'd91509: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=92;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=1134;
 end   
19'd91510: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=9;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=2643;
 end   
19'd91511: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd91512: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=76;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16963;
 end   
19'd91513: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=92;
   mapp<=71;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=13496;
 end   
19'd91514: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=80;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=17425;
 end   
19'd91515: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=64;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=10726;
 end   
19'd91516: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=41;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=6597;
 end   
19'd91517: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=26;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=10800;
 end   
19'd91518: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=86;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=10140;
 end   
19'd91519: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=35;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=11858;
 end   
19'd91520: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=33;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=8334;
 end   
19'd91521: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=51;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=8727;
 end   
19'd91522: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd91523: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd91665: begin  
rid<=1;
end
19'd91666: begin  
end
19'd91667: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd91668: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd91669: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd91670: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd91671: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd91672: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd91673: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd91674: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd91675: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd91676: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd91677: begin  
rid<=0;
end
19'd91801: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=10;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13093;
 end   
19'd91802: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=83;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd91803: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=3;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd91804: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=37;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd91805: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=83;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd91806: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=41;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd91807: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=35;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd91808: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=21;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd91809: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=77;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd91810: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=48;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=28544;
 end   
19'd91811: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=32;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd91812: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=41;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd91813: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=70;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd91814: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=16;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd91815: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=63;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd91816: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=18;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd91817: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=15;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd91818: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=84;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd91819: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd91961: begin  
rid<=1;
end
19'd91962: begin  
end
19'd91963: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd91964: begin  
rid<=0;
end
19'd92101: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=96;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3936;
 end   
19'd92102: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=85;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8170;
 end   
19'd92103: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=8;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=788;
 end   
19'd92104: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=60;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5790;
 end   
19'd92105: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=48;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4648;
 end   
19'd92106: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=85;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=8210;
 end   
19'd92107: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=78;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=7548;
 end   
19'd92108: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=1;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=166;
 end   
19'd92109: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=71;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=6896;
 end   
19'd92110: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=5;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=570;
 end   
19'd92111: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=1;
   pp<=100;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[10]<=196;
 end   
19'd92112: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=52;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7680;
 end   
19'd92113: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=9;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8638;
 end   
19'd92114: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=31;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=2400;
 end   
19'd92115: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=87;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=10314;
 end   
19'd92116: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=70;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=8288;
 end   
19'd92117: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=25;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=9510;
 end   
19'd92118: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=84;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=11916;
 end   
19'd92119: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=2;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=270;
 end   
19'd92120: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=27;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=8300;
 end   
19'd92121: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=46;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=2962;
 end   
19'd92122: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=88;
   pp<=100;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[10]<=4772;
 end   
19'd92123: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd92265: begin  
rid<=1;
end
19'd92266: begin  
end
19'd92267: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd92268: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd92269: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd92270: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd92271: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd92272: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd92273: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd92274: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd92275: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd92276: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd92277: begin  
check0<=expctdoutput[10]-outcheck0;
end
19'd92278: begin  
rid<=0;
end
19'd92401: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=51;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6609;
 end   
19'd92402: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=18;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd92403: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=19;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12157;
 end   
19'd92404: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=73;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd92405: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd92547: begin  
rid<=1;
end
19'd92548: begin  
end
19'd92549: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd92550: begin  
rid<=0;
end
19'd92701: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=59;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16835;
 end   
19'd92702: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=18;
   mapp<=10;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=17792;
 end   
19'd92703: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=61;
   mapp<=59;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=21437;
 end   
19'd92704: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=67;
   mapp<=25;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=24762;
 end   
19'd92705: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=3;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd92706: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=66;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd92707: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=38;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd92708: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=26;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd92709: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=93;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd92710: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=82;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd92711: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=76;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd92712: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=21;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=38442;
 end   
19'd92713: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=73;
   mapp<=38;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=44434;
 end   
19'd92714: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=98;
   mapp<=57;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=43334;
 end   
19'd92715: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=57;
   mapp<=80;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=46849;
 end   
19'd92716: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=58;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd92717: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=19;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd92718: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=45;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd92719: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=1;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd92720: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd92721: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd92722: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=56;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd92723: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd92865: begin  
rid<=1;
end
19'd92866: begin  
end
19'd92867: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd92868: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd92869: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd92870: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd92871: begin  
rid<=0;
end
19'd93001: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=38;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11085;
 end   
19'd93002: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=30;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=16272;
 end   
19'd93003: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=5;
   mapp<=78;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=17173;
 end   
19'd93004: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=90;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd93005: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=99;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd93006: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=69;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd93007: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=7;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd93008: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=53;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd93009: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=13;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd93010: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=56;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd93011: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=35;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=36500;
 end   
19'd93012: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=19;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=40773;
 end   
19'd93013: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=71;
   mapp<=48;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=40413;
 end   
19'd93014: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=64;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd93015: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=99;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd93016: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=8;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd93017: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=47;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd93018: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=14;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd93019: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=14;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd93020: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd93021: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd93163: begin  
rid<=1;
end
19'd93164: begin  
end
19'd93165: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd93166: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd93167: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd93168: begin  
rid<=0;
end
19'd93301: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=86;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=22109;
 end   
19'd93302: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=92;
   mapp<=92;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=25221;
 end   
19'd93303: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=52;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd93304: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=17;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd93305: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=24;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd93306: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=88;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd93307: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=93;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd93308: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=58;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=45431;
 end   
19'd93309: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=37;
   mapp<=88;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=46600;
 end   
19'd93310: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=45;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd93311: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=68;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd93312: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=97;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd93313: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=25;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd93314: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=47;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd93315: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd93457: begin  
rid<=1;
end
19'd93458: begin  
end
19'd93459: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd93460: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd93461: begin  
rid<=0;
end
19'd93601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=12;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14051;
 end   
19'd93602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=20;
   mapp<=7;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=18919;
 end   
19'd93603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=31;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=16243;
 end   
19'd93604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=76;
   mapp<=49;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=16916;
 end   
19'd93605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=91;
   mapp<=46;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=18663;
 end   
19'd93606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=25;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd93607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=45;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd93608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=99;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd93609: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd93610: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=74;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd93611: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=56;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd93612: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=58;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=31160;
 end   
19'd93613: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=88;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=32888;
 end   
19'd93614: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=44;
   mapp<=36;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=28266;
 end   
19'd93615: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=4;
   mapp<=8;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=25552;
 end   
19'd93616: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=30;
   mapp<=96;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=32059;
 end   
19'd93617: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=27;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd93618: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=49;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd93619: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=19;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd93620: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=68;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd93621: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=74;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd93622: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=1;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd93623: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd93765: begin  
rid<=1;
end
19'd93766: begin  
end
19'd93767: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd93768: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd93769: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd93770: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd93771: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd93772: begin  
rid<=0;
end
19'd93901: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=13;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2532;
 end   
19'd93902: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=62;
   mapp<=27;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6262;
 end   
19'd93903: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=80;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5786;
 end   
19'd93904: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=18;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1974;
 end   
19'd93905: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=28;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4291;
 end   
19'd93906: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=89;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6275;
 end   
19'd93907: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=13;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=2025;
 end   
19'd93908: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=41;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=3397;
 end   
19'd93909: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=23;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=4190;
 end   
19'd93910: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=96;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd93911: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=31;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=4893;
 end   
19'd93912: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=35;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8627;
 end   
19'd93913: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=32;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=10058;
 end   
19'd93914: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=82;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=7796;
 end   
19'd93915: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=82;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=8833;
 end   
19'd93916: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=50;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=9585;
 end   
19'd93917: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=44;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=5469;
 end   
19'd93918: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=52;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=7289;
 end   
19'd93919: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=57;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=5997;
 end   
19'd93920: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=1;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd93921: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd94063: begin  
rid<=1;
end
19'd94064: begin  
end
19'd94065: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd94066: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd94067: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd94068: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd94069: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd94070: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd94071: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd94072: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd94073: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd94074: begin  
rid<=0;
end
19'd94201: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=82;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7114;
 end   
19'd94202: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=12;
   mapp<=94;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7946;
 end   
19'd94203: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=19;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1890;
 end   
19'd94204: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=26;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3158;
 end   
19'd94205: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=83;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=7242;
 end   
19'd94206: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd94207: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=96;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=10620;
 end   
19'd94208: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=2;
   mapp<=25;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=10450;
 end   
19'd94209: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=52;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=6906;
 end   
19'd94210: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=12;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=4358;
 end   
19'd94211: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=24;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=9636;
 end   
19'd94212: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd94213: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd94355: begin  
rid<=1;
end
19'd94356: begin  
end
19'd94357: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd94358: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd94359: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd94360: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd94361: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd94362: begin  
rid<=0;
end
19'd94501: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=11;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9192;
 end   
19'd94502: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=81;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8325;
 end   
19'd94503: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=50;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd94504: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd94505: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=59;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17379;
 end   
19'd94506: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=16;
   mapp<=53;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=15232;
 end   
19'd94507: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=97;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd94508: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=18;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd94509: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd94651: begin  
rid<=1;
end
19'd94652: begin  
end
19'd94653: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd94654: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd94655: begin  
rid<=0;
end
19'd94801: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=41;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13164;
 end   
19'd94802: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=9;
   mapp<=65;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12454;
 end   
19'd94803: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=97;
   mapp<=52;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=17996;
 end   
19'd94804: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=62;
   mapp<=13;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=17458;
 end   
19'd94805: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=48;
   mapp<=71;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=18581;
 end   
19'd94806: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd94807: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd94808: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd94809: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd94810: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=38;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=23400;
 end   
19'd94811: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=6;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18825;
 end   
19'd94812: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=61;
   mapp<=92;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=25141;
 end   
19'd94813: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=50;
   mapp<=36;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=22561;
 end   
19'd94814: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=47;
   mapp<=20;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=26219;
 end   
19'd94815: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd94816: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd94817: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd94818: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd94819: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd94961: begin  
rid<=1;
end
19'd94962: begin  
end
19'd94963: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd94964: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd94965: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd94966: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd94967: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd94968: begin  
rid<=0;
end
19'd95101: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=1;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8631;
 end   
19'd95102: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=16;
   mapp<=81;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12890;
 end   
19'd95103: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=94;
   mapp<=68;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9915;
 end   
19'd95104: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=67;
   mapp<=14;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=9112;
 end   
19'd95105: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=45;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=9226;
 end   
19'd95106: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=67;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7828;
 end   
19'd95107: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=39;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=6394;
 end   
19'd95108: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=63;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd95109: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd95110: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=74;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd95111: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=17;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=19860;
 end   
19'd95112: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=24;
   mapp<=99;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=26867;
 end   
19'd95113: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=49;
   mapp<=25;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=26995;
 end   
19'd95114: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=86;
   mapp<=80;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=28447;
 end   
19'd95115: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=74;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=21450;
 end   
19'd95116: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=57;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=23766;
 end   
19'd95117: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=85;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=19069;
 end   
19'd95118: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=15;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd95119: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=58;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd95120: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=75;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd95121: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd95263: begin  
rid<=1;
end
19'd95264: begin  
end
19'd95265: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd95266: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd95267: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd95268: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd95269: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd95270: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd95271: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd95272: begin  
rid<=0;
end
19'd95401: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=61;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12547;
 end   
19'd95402: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=12;
   mapp<=37;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15975;
 end   
19'd95403: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=96;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd95404: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=76;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd95405: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd95406: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd95407: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=50;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=25197;
 end   
19'd95408: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=58;
   mapp<=71;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=31253;
 end   
19'd95409: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=28;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd95410: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=45;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd95411: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=42;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd95412: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd95413: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd95555: begin  
rid<=1;
end
19'd95556: begin  
end
19'd95557: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd95558: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd95559: begin  
rid<=0;
end
19'd95701: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=95;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8452;
 end   
19'd95702: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=4;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd95703: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=13;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd95704: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=95;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12209;
 end   
19'd95705: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=21;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd95706: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=48;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd95707: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd95849: begin  
rid<=1;
end
19'd95850: begin  
end
19'd95851: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd95852: begin  
rid<=0;
end
19'd96001: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=19;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3747;
 end   
19'd96002: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=37;
   mapp<=91;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3145;
 end   
19'd96003: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=38;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1926;
 end   
19'd96004: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd96005: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=31;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=6977;
 end   
19'd96006: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=37;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=6431;
 end   
19'd96007: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=62;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=5106;
 end   
19'd96008: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd96009: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd96151: begin  
rid<=1;
end
19'd96152: begin  
end
19'd96153: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd96154: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd96155: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd96156: begin  
rid<=0;
end
19'd96301: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=11;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11262;
 end   
19'd96302: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=97;
   mapp<=14;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10796;
 end   
19'd96303: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=37;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd96304: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=2;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd96305: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=15;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd96306: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=63;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd96307: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=17;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd96308: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=17;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd96309: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=99;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd96310: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd96311: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=74;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=31324;
 end   
19'd96312: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=91;
   mapp<=43;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=26252;
 end   
19'd96313: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=8;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd96314: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=18;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd96315: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=51;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd96316: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=77;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd96317: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=23;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd96318: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=52;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd96319: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=11;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd96320: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd96321: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd96463: begin  
rid<=1;
end
19'd96464: begin  
end
19'd96465: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd96466: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd96467: begin  
rid<=0;
end
19'd96601: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=21;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1326;
 end   
19'd96602: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=87;
   mapp<=15;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7894;
 end   
19'd96603: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=87;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4283;
 end   
19'd96604: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=28;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3141;
 end   
19'd96605: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd96606: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=46;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=6249;
 end   
19'd96607: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=75;
   mapp<=27;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=15736;
 end   
19'd96608: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=88;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=14106;
 end   
19'd96609: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=77;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=7733;
 end   
19'd96610: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd96611: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd96753: begin  
rid<=1;
end
19'd96754: begin  
end
19'd96755: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd96756: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd96757: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd96758: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd96759: begin  
rid<=0;
end
19'd96901: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=69;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3584;
 end   
19'd96902: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=47;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd96903: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=60;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7616;
 end   
19'd96904: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=52;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd96905: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd97047: begin  
rid<=1;
end
19'd97048: begin  
end
19'd97049: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd97050: begin  
rid<=0;
end
19'd97201: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=51;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11697;
 end   
19'd97202: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=5;
   mapp<=80;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12831;
 end   
19'd97203: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=40;
   mapp<=41;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=17155;
 end   
19'd97204: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=89;
   mapp<=50;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=13199;
 end   
19'd97205: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=25;
   mapp<=39;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=14438;
 end   
19'd97206: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=82;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd97207: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=4;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd97208: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=53;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd97209: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=80;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd97210: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=30;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd97211: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=11;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd97212: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=47;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=23188;
 end   
19'd97213: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=7;
   mapp<=58;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=21637;
 end   
19'd97214: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=96;
   mapp<=87;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=22269;
 end   
19'd97215: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=14;
   mapp<=51;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=19632;
 end   
19'd97216: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=5;
   mapp<=27;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=21733;
 end   
19'd97217: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=49;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd97218: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=6;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd97219: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=10;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd97220: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=15;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd97221: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=35;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd97222: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd97223: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd97365: begin  
rid<=1;
end
19'd97366: begin  
end
19'd97367: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd97368: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd97369: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd97370: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd97371: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd97372: begin  
rid<=0;
end
19'd97501: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=66;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10461;
 end   
19'd97502: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=27;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd97503: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=25;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd97504: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd97505: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=48;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd97506: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=75;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd97507: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=30;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd97508: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=57;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd97509: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=13;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd97510: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=52;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=34369;
 end   
19'd97511: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=55;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd97512: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=84;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd97513: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=35;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd97514: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=94;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd97515: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=46;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd97516: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=90;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd97517: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=36;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd97518: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=47;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd97519: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd97661: begin  
rid<=1;
end
19'd97662: begin  
end
19'd97663: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd97664: begin  
rid<=0;
end
19'd97801: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=46;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11112;
 end   
19'd97802: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=99;
   mapp<=58;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=16460;
 end   
19'd97803: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=22;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd97804: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=92;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd97805: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=41;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16325;
 end   
19'd97806: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=91;
   mapp<=8;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=19499;
 end   
19'd97807: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=76;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd97808: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=24;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd97809: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd97951: begin  
rid<=1;
end
19'd97952: begin  
end
19'd97953: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd97954: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd97955: begin  
rid<=0;
end
19'd98101: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=37;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=20363;
 end   
19'd98102: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=9;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd98103: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=50;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd98104: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=54;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd98105: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=40;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd98106: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=97;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd98107: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=27;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd98108: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=79;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd98109: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=46;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd98110: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=39;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd98111: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=93;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=57922;
 end   
19'd98112: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=51;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd98113: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=16;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd98114: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=94;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd98115: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=38;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd98116: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=88;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd98117: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=75;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd98118: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=71;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd98119: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=21;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd98120: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=80;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd98121: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd98263: begin  
rid<=1;
end
19'd98264: begin  
end
19'd98265: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd98266: begin  
rid<=0;
end
19'd98401: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=56;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5544;
 end   
19'd98402: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=9;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=901;
 end   
19'd98403: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=66;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6554;
 end   
19'd98404: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=68;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6762;
 end   
19'd98405: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=59;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5881;
 end   
19'd98406: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=95;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=9455;
 end   
19'd98407: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=28;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7896;
 end   
19'd98408: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=94;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8797;
 end   
19'd98409: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=32;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=9242;
 end   
19'd98410: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=66;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=12306;
 end   
19'd98411: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=58;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=10753;
 end   
19'd98412: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=66;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=14999;
 end   
19'd98413: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd98555: begin  
rid<=1;
end
19'd98556: begin  
end
19'd98557: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd98558: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd98559: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd98560: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd98561: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd98562: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd98563: begin  
rid<=0;
end
19'd98701: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=49;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12489;
 end   
19'd98702: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=22;
   mapp<=86;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15650;
 end   
19'd98703: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=60;
   mapp<=60;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=17754;
 end   
19'd98704: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=83;
   mapp<=66;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=13237;
 end   
19'd98705: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=73;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=11375;
 end   
19'd98706: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=66;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd98707: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=6;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd98708: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=46;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd98709: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=20;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=23131;
 end   
19'd98710: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=66;
   mapp<=8;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=26564;
 end   
19'd98711: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=69;
   mapp<=46;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=27386;
 end   
19'd98712: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=78;
   mapp<=70;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=26853;
 end   
19'd98713: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=27;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=21671;
 end   
19'd98714: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd98715: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=84;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd98716: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=59;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd98717: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd98859: begin  
rid<=1;
end
19'd98860: begin  
end
19'd98861: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd98862: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd98863: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd98864: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd98865: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd98866: begin  
rid<=0;
end
19'd99001: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=93;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5163;
 end   
19'd99002: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=44;
   mapp<=21;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5756;
 end   
19'd99003: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=9;
   mapp<=91;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6147;
 end   
19'd99004: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=7;
   mapp<=90;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5153;
 end   
19'd99005: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=40;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=7955;
 end   
19'd99006: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=23;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=9979;
 end   
19'd99007: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=22;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=8507;
 end   
19'd99008: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=47;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=10385;
 end   
19'd99009: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=50;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd99010: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=25;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd99011: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd99012: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=55;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=11145;
 end   
19'd99013: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=5;
   mapp<=69;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=11503;
 end   
19'd99014: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=26;
   mapp<=40;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=16881;
 end   
19'd99015: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=87;
   mapp<=1;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=19860;
 end   
19'd99016: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=63;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=21290;
 end   
19'd99017: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=79;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=24176;
 end   
19'd99018: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=66;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=21110;
 end   
19'd99019: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=78;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=20332;
 end   
19'd99020: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=45;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd99021: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=9;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd99022: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=86;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd99023: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd99165: begin  
rid<=1;
end
19'd99166: begin  
end
19'd99167: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd99168: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd99169: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd99170: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd99171: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd99172: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd99173: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd99174: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd99175: begin  
rid<=0;
end
19'd99301: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=61;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4717;
 end   
19'd99302: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=83;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd99303: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=38;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd99304: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=99;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16470;
 end   
19'd99305: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=97;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd99306: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=95;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd99307: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd99449: begin  
rid<=1;
end
19'd99450: begin  
end
19'd99451: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd99452: begin  
rid<=0;
end
19'd99601: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=89;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5963;
 end   
19'd99602: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3570;
 end   
19'd99603: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=3;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=287;
 end   
19'd99604: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=55;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4925;
 end   
19'd99605: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=55;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4935;
 end   
19'd99606: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=52;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=4678;
 end   
19'd99607: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=56;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=5044;
 end   
19'd99608: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=45;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=4075;
 end   
19'd99609: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=62;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=5598;
 end   
19'd99610: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=97;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=8723;
 end   
19'd99611: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=50;
   pp<=100;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[10]<=4550;
 end   
19'd99612: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=3;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=6158;
 end   
19'd99613: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=3585;
 end   
19'd99614: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=27;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=368;
 end   
19'd99615: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=47;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=5066;
 end   
19'd99616: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=27;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=5016;
 end   
19'd99617: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=3;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=4687;
 end   
19'd99618: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=76;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=5272;
 end   
19'd99619: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=65;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=4270;
 end   
19'd99620: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=75;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=5823;
 end   
19'd99621: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=46;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=8861;
 end   
19'd99622: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=81;
   pp<=100;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[10]<=4793;
 end   
19'd99623: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd99765: begin  
rid<=1;
end
19'd99766: begin  
end
19'd99767: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd99768: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd99769: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd99770: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd99771: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd99772: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd99773: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd99774: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd99775: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd99776: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd99777: begin  
check0<=expctdoutput[10]-outcheck0;
end
19'd99778: begin  
rid<=0;
end
19'd99901: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=74;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=18243;
 end   
19'd99902: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=8;
   mapp<=16;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=14897;
 end   
19'd99903: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=35;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd99904: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=2;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd99905: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=35;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd99906: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=41;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd99907: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=86;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd99908: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=93;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd99909: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=20;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd99910: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd99911: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=83;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=30258;
 end   
19'd99912: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=33;
   mapp<=44;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=30133;
 end   
19'd99913: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=11;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd99914: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=76;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd99915: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=5;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd99916: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=65;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd99917: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=6;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd99918: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=98;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd99919: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=18;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd99920: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd99921: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd100063: begin  
rid<=1;
end
19'd100064: begin  
end
19'd100065: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd100066: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd100067: begin  
rid<=0;
end
19'd100201: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=65;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=19786;
 end   
19'd100202: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=62;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=20201;
 end   
19'd100203: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=39;
   mapp<=50;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=21891;
 end   
19'd100204: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=8;
   mapp<=34;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=24429;
 end   
19'd100205: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=60;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd100206: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=82;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd100207: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd100208: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd100209: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd100210: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=73;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=40865;
 end   
19'd100211: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=50;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=38703;
 end   
19'd100212: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=60;
   mapp<=22;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=34137;
 end   
19'd100213: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=41;
   mapp<=35;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=40405;
 end   
19'd100214: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=93;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd100215: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=48;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd100216: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd100217: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd100218: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd100219: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd100361: begin  
rid<=1;
end
19'd100362: begin  
end
19'd100363: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd100364: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd100365: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd100366: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd100367: begin  
rid<=0;
end
19'd100501: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=12;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=816;
 end   
19'd100502: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=65;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4430;
 end   
19'd100503: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=19;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1312;
 end   
19'd100504: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=27;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1866;
 end   
19'd100505: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=71;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4868;
 end   
19'd100506: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=14;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=1002;
 end   
19'd100507: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=42;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=2916;
 end   
19'd100508: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=50;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=3470;
 end   
19'd100509: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=28;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=2188;
 end   
19'd100510: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=61;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=7419;
 end   
19'd100511: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=77;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=5085;
 end   
19'd100512: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=36;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=3630;
 end   
19'd100513: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=25;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=6093;
 end   
19'd100514: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=6;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=1296;
 end   
19'd100515: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=65;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=6101;
 end   
19'd100516: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=83;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=7537;
 end   
19'd100517: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd100659: begin  
rid<=1;
end
19'd100660: begin  
end
19'd100661: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd100662: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd100663: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd100664: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd100665: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd100666: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd100667: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd100668: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd100669: begin  
rid<=0;
end
19'd100801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=31;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=19657;
 end   
19'd100802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=80;
   mapp<=53;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=17806;
 end   
19'd100803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=83;
   mapp<=65;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=15030;
 end   
19'd100804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=47;
   mapp<=45;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=15679;
 end   
19'd100805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=23;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd100806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=81;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd100807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=63;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd100808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=44;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd100809: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=49;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd100810: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=98;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=37776;
 end   
19'd100811: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=78;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=37765;
 end   
19'd100812: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=27;
   mapp<=62;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=31305;
 end   
19'd100813: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=25;
   mapp<=91;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=35560;
 end   
19'd100814: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=60;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd100815: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=69;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd100816: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=80;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd100817: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd100818: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=47;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd100819: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd100961: begin  
rid<=1;
end
19'd100962: begin  
end
19'd100963: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd100964: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd100965: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd100966: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd100967: begin  
rid<=0;
end
19'd101101: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=23;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1886;
 end   
19'd101102: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=87;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=6671;
 end   
19'd101103: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd101245: begin  
rid<=1;
end
19'd101246: begin  
end
19'd101247: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd101248: begin  
rid<=0;
end
19'd101401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=56;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=20497;
 end   
19'd101402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=24;
   mapp<=91;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=18535;
 end   
19'd101403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=17;
   mapp<=11;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=24226;
 end   
19'd101404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=56;
   mapp<=44;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=25267;
 end   
19'd101405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=48;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd101406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=60;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd101407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=80;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd101408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=50;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd101409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd101410: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=66;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd101411: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=67;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd101412: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=35;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=46401;
 end   
19'd101413: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=16;
   mapp<=73;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=44341;
 end   
19'd101414: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=57;
   mapp<=43;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=55855;
 end   
19'd101415: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=80;
   mapp<=48;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=56831;
 end   
19'd101416: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=66;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd101417: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=61;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd101418: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=91;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd101419: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=33;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd101420: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=29;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd101421: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=85;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd101422: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=50;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd101423: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd101565: begin  
rid<=1;
end
19'd101566: begin  
end
19'd101567: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd101568: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd101569: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd101570: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd101571: begin  
rid<=0;
end
19'd101701: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=88;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7744;
 end   
19'd101702: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=86;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7578;
 end   
19'd101703: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=57;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5036;
 end   
19'd101704: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=59;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5222;
 end   
19'd101705: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=27;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2416;
 end   
19'd101706: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=10;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=930;
 end   
19'd101707: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=26;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=2348;
 end   
19'd101708: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=90;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=7990;
 end   
19'd101709: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=64;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=10368;
 end   
19'd101710: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=66;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=10284;
 end   
19'd101711: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=74;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=8070;
 end   
19'd101712: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=92;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=8994;
 end   
19'd101713: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=48;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=4384;
 end   
19'd101714: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=12;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=1422;
 end   
19'd101715: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=92;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=6120;
 end   
19'd101716: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=16;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=8646;
 end   
19'd101717: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd101859: begin  
rid<=1;
end
19'd101860: begin  
end
19'd101861: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd101862: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd101863: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd101864: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd101865: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd101866: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd101867: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd101868: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd101869: begin  
rid<=0;
end
19'd102001: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=96;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=21072;
 end   
19'd102002: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=96;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd102003: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=78;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd102004: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=8;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd102005: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=86;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd102006: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=37;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd102007: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=3;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd102008: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=93;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=30815;
 end   
19'd102009: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=54;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd102010: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=94;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd102011: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=4;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd102012: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=42;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd102013: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=24;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd102014: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=69;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd102015: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd102157: begin  
rid<=1;
end
19'd102158: begin  
end
19'd102159: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd102160: begin  
rid<=0;
end
19'd102301: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=2;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=77;
 end   
19'd102302: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=23;
   mapp<=1;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=669;
 end   
19'd102303: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=38;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1107;
 end   
19'd102304: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=61;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd102305: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=5;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=247;
 end   
19'd102306: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=0;
   mapp<=1;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=701;
 end   
19'd102307: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=32;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=2251;
 end   
19'd102308: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=56;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd102309: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd102451: begin  
rid<=1;
end
19'd102452: begin  
end
19'd102453: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd102454: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd102455: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd102456: begin  
rid<=0;
end
19'd102601: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=92;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2494;
 end   
19'd102602: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=10;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9336;
 end   
19'd102603: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd102604: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=89;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=11056;
 end   
19'd102605: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=69;
   mapp<=8;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=15223;
 end   
19'd102606: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd102607: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd102749: begin  
rid<=1;
end
19'd102750: begin  
end
19'd102751: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd102752: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd102753: begin  
rid<=0;
end
19'd102901: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=36;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1908;
 end   
19'd102902: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=95;
   mapp<=6;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4077;
 end   
19'd102903: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=2;
   mapp<=39;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8497;
 end   
19'd102904: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=73;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=9359;
 end   
19'd102905: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=69;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=9547;
 end   
19'd102906: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=73;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6912;
 end   
19'd102907: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=44;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=4399;
 end   
19'd102908: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd102909: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd102910: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=57;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=3831;
 end   
19'd102911: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=47;
   mapp<=7;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=7494;
 end   
19'd102912: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=31;
   mapp<=22;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=14247;
 end   
19'd102913: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=64;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=15511;
 end   
19'd102914: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=48;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=14891;
 end   
19'd102915: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=8;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=11000;
 end   
19'd102916: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=72;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=11669;
 end   
19'd102917: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd102918: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd102919: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd103061: begin  
rid<=1;
end
19'd103062: begin  
end
19'd103063: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd103064: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd103065: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd103066: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd103067: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd103068: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd103069: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd103070: begin  
rid<=0;
end
19'd103201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=90;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5099;
 end   
19'd103202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=67;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=901;
 end   
19'd103203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=5;
   mapp<=14;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1949;
 end   
19'd103204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=11;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6399;
 end   
19'd103205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=83;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd103206: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=53;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd103207: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=29;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8404;
 end   
19'd103208: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=40;
   mapp<=26;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=4843;
 end   
19'd103209: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=27;
   mapp<=42;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=7654;
 end   
19'd103210: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=40;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=12001;
 end   
19'd103211: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=86;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd103212: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=43;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd103213: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd103355: begin  
rid<=1;
end
19'd103356: begin  
end
19'd103357: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd103358: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd103359: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd103360: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd103361: begin  
rid<=0;
end
19'd103501: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=42;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11176;
 end   
19'd103502: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=32;
   mapp<=10;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10024;
 end   
19'd103503: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=42;
   mapp<=5;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11540;
 end   
19'd103504: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=20;
   mapp<=9;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=12116;
 end   
19'd103505: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=25;
   mapp<=71;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=10795;
 end   
19'd103506: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=81;
   mapp<=71;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=14538;
 end   
19'd103507: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=18;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd103508: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd103509: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=51;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd103510: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=52;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd103511: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=57;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd103512: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=88;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=28059;
 end   
19'd103513: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=47;
   mapp<=75;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=26832;
 end   
19'd103514: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=72;
   mapp<=30;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=27593;
 end   
19'd103515: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=90;
   mapp<=51;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=27564;
 end   
19'd103516: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=19;
   mapp<=2;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=23867;
 end   
19'd103517: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=17;
   mapp<=50;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=32108;
 end   
19'd103518: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=93;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd103519: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=60;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd103520: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=56;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd103521: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=92;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd103522: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=93;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd103523: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd103665: begin  
rid<=1;
end
19'd103666: begin  
end
19'd103667: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd103668: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd103669: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd103670: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd103671: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd103672: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd103673: begin  
rid<=0;
end
19'd103801: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=44;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10767;
 end   
19'd103802: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=56;
   mapp<=73;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12219;
 end   
19'd103803: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=86;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd103804: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=25;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd103805: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=64;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd103806: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=53;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=15260;
 end   
19'd103807: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=9;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=16653;
 end   
19'd103808: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=95;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd103809: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=47;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd103810: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=8;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd103811: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd103953: begin  
rid<=1;
end
19'd103954: begin  
end
19'd103955: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd103956: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd103957: begin  
rid<=0;
end
19'd104101: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=82;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8322;
 end   
19'd104102: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=90;
   mapp<=23;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6999;
 end   
19'd104103: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=75;
   mapp<=44;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5494;
 end   
19'd104104: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=46;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4695;
 end   
19'd104105: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=39;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5408;
 end   
19'd104106: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=48;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6001;
 end   
19'd104107: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=65;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=6818;
 end   
19'd104108: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=62;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=4702;
 end   
19'd104109: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=68;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd104110: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=19;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd104111: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=87;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=18463;
 end   
19'd104112: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=40;
   mapp<=82;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=15600;
 end   
19'd104113: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=66;
   mapp<=13;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=13924;
 end   
19'd104114: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=33;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=14625;
 end   
19'd104115: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=90;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=13808;
 end   
19'd104116: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=21;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=11403;
 end   
19'd104117: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=36;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=16851;
 end   
19'd104118: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=77;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=17883;
 end   
19'd104119: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=95;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd104120: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=6;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd104121: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd104263: begin  
rid<=1;
end
19'd104264: begin  
end
19'd104265: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd104266: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd104267: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd104268: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd104269: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd104270: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd104271: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd104272: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd104273: begin  
rid<=0;
end
19'd104401: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=57;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4329;
 end   
19'd104402: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=21;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7921;
 end   
19'd104403: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=61;
   mapp<=33;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6642;
 end   
19'd104404: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd104405: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd104406: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=78;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=10771;
 end   
19'd104407: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=97;
   mapp<=60;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=16295;
 end   
19'd104408: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=34;
   mapp<=16;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15293;
 end   
19'd104409: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd104410: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd104411: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd104553: begin  
rid<=1;
end
19'd104554: begin  
end
19'd104555: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd104556: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd104557: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd104558: begin  
rid<=0;
end
19'd104701: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=37;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=24820;
 end   
19'd104702: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=99;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=26650;
 end   
19'd104703: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=48;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd104704: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=93;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd104705: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=58;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd104706: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=57;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd104707: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=71;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd104708: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=58;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd104709: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=82;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd104710: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=36;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=37162;
 end   
19'd104711: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=43;
   mapp<=65;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=35323;
 end   
19'd104712: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=16;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd104713: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=78;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd104714: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=6;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd104715: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=24;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd104716: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=15;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd104717: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=73;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd104718: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=60;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd104719: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd104861: begin  
rid<=1;
end
19'd104862: begin  
end
19'd104863: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd104864: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd104865: begin  
rid<=0;
end
19'd105001: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=21;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3535;
 end   
19'd105002: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=16;
   mapp<=8;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8606;
 end   
19'd105003: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=23;
   mapp<=88;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=13861;
 end   
19'd105004: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=12;
   mapp<=82;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=12518;
 end   
19'd105005: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=86;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd105006: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd105007: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=66;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd105008: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=62;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17993;
 end   
19'd105009: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=46;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=19424;
 end   
19'd105010: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=81;
   mapp<=58;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=23987;
 end   
19'd105011: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=53;
   mapp<=76;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=24592;
 end   
19'd105012: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=4;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd105013: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd105014: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=97;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd105015: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd105157: begin  
rid<=1;
end
19'd105158: begin  
end
19'd105159: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd105160: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd105161: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd105162: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd105163: begin  
rid<=0;
end
19'd105301: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=31;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10357;
 end   
19'd105302: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=65;
   mapp<=15;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10674;
 end   
19'd105303: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=56;
   mapp<=87;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11560;
 end   
19'd105304: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=84;
   mapp<=21;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=12462;
 end   
19'd105305: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=65;
   mapp<=37;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=13335;
 end   
19'd105306: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=4;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=17150;
 end   
19'd105307: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=78;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=20316;
 end   
19'd105308: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd105309: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd105310: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd105311: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd105312: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=86;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17435;
 end   
19'd105313: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=43;
   mapp<=65;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20334;
 end   
19'd105314: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=35;
   mapp<=0;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=18652;
 end   
19'd105315: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=12;
   mapp<=84;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=25482;
 end   
19'd105316: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=31;
   mapp<=89;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=22361;
 end   
19'd105317: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=2;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=20091;
 end   
19'd105318: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=11;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=24879;
 end   
19'd105319: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd105320: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd105321: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd105322: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd105323: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd105465: begin  
rid<=1;
end
19'd105466: begin  
end
19'd105467: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd105468: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd105469: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd105470: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd105471: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd105472: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd105473: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd105474: begin  
rid<=0;
end
19'd105601: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=90;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12651;
 end   
19'd105602: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=64;
   mapp<=1;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9324;
 end   
19'd105603: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=97;
   mapp<=35;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=13101;
 end   
19'd105604: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=25;
   mapp<=46;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=16789;
 end   
19'd105605: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=7;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd105606: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=83;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd105607: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=15;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd105608: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=77;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd105609: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=94;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd105610: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=80;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd105611: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=55;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd105612: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=41;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=26415;
 end   
19'd105613: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=60;
   mapp<=34;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=23531;
 end   
19'd105614: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=73;
   mapp<=83;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=30959;
 end   
19'd105615: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=23;
   mapp<=11;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=27786;
 end   
19'd105616: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=89;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd105617: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=32;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd105618: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=23;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd105619: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=87;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd105620: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=78;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd105621: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=39;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd105622: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=3;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd105623: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd105765: begin  
rid<=1;
end
19'd105766: begin  
end
19'd105767: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd105768: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd105769: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd105770: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd105771: begin  
rid<=0;
end
19'd105901: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=14;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10396;
 end   
19'd105902: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=99;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=17011;
 end   
19'd105903: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=98;
   mapp<=1;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9784;
 end   
19'd105904: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=3;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd105905: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=98;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd105906: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=17;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd105907: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=90;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd105908: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=68;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd105909: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=26;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=30082;
 end   
19'd105910: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=67;
   mapp<=92;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=32191;
 end   
19'd105911: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=35;
   mapp<=48;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=19000;
 end   
19'd105912: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=7;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd105913: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=77;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd105914: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=71;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd105915: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=5;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd105916: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=30;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd105917: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd106059: begin  
rid<=1;
end
19'd106060: begin  
end
19'd106061: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd106062: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd106063: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd106064: begin  
rid<=0;
end
19'd106201: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=59;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3422;
 end   
19'd106202: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=98;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5694;
 end   
19'd106203: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=42;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2456;
 end   
19'd106204: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=8;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=494;
 end   
19'd106205: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=77;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4506;
 end   
19'd106206: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=33;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5600;
 end   
19'd106207: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=5;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=6024;
 end   
19'd106208: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=78;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=7604;
 end   
19'd106209: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=90;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6434;
 end   
19'd106210: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=11;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=5232;
 end   
19'd106211: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd106353: begin  
rid<=1;
end
19'd106354: begin  
end
19'd106355: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd106356: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd106357: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd106358: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd106359: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd106360: begin  
rid<=0;
end
19'd106501: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=60;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11310;
 end   
19'd106502: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=57;
   mapp<=69;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12537;
 end   
19'd106503: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=63;
   mapp<=43;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11130;
 end   
19'd106504: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=46;
   mapp<=48;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=12740;
 end   
19'd106505: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=90;
   mapp<=26;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=10418;
 end   
19'd106506: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=68;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd106507: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=26;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd106508: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=86;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd106509: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=10;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd106510: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=20;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=22754;
 end   
19'd106511: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=37;
   mapp<=39;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=24782;
 end   
19'd106512: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=15;
   mapp<=13;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=25658;
 end   
19'd106513: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=75;
   mapp<=62;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=27473;
 end   
19'd106514: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=72;
   mapp<=58;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=23068;
 end   
19'd106515: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=76;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd106516: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=90;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd106517: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=29;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd106518: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=55;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd106519: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd106661: begin  
rid<=1;
end
19'd106662: begin  
end
19'd106663: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd106664: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd106665: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd106666: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd106667: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd106668: begin  
rid<=0;
end
19'd106801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=90;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=15192;
 end   
19'd106802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=33;
   mapp<=75;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=14487;
 end   
19'd106803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=67;
   mapp<=35;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10134;
 end   
19'd106804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=37;
   mapp<=76;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=12479;
 end   
19'd106805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd106806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd106807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd106808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=75;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=18931;
 end   
19'd106809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=41;
   mapp<=45;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20421;
 end   
19'd106810: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=25;
   mapp<=3;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=16397;
 end   
19'd106811: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=1;
   mapp<=94;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=23957;
 end   
19'd106812: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd106813: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd106814: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd106815: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd106957: begin  
rid<=1;
end
19'd106958: begin  
end
19'd106959: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd106960: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd106961: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd106962: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd106963: begin  
rid<=0;
end
19'd107101: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=26;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12613;
 end   
19'd107102: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=25;
   mapp<=91;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10826;
 end   
19'd107103: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=90;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd107104: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=89;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd107105: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=0;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd107106: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=14;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=15214;
 end   
19'd107107: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=28;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=16863;
 end   
19'd107108: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=13;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd107109: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=48;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd107110: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=0;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd107111: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd107253: begin  
rid<=1;
end
19'd107254: begin  
end
19'd107255: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd107256: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd107257: begin  
rid<=0;
end
19'd107401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=50;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5325;
 end   
19'd107402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=53;
   mapp<=9;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7403;
 end   
19'd107403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=53;
   mapp<=66;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10210;
 end   
19'd107404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=65;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=11336;
 end   
19'd107405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=65;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=11770;
 end   
19'd107406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=87;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=12297;
 end   
19'd107407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd107408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd107409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=88;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8575;
 end   
19'd107410: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=68;
   mapp<=9;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=11119;
 end   
19'd107411: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=2;
   mapp<=43;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=14136;
 end   
19'd107412: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=16186;
 end   
19'd107413: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=71;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=18922;
 end   
19'd107414: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=11;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=18695;
 end   
19'd107415: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd107416: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd107417: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd107559: begin  
rid<=1;
end
19'd107560: begin  
end
19'd107561: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd107562: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd107563: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd107564: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd107565: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd107566: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd107567: begin  
rid<=0;
end
19'd107701: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=13;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14676;
 end   
19'd107702: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=96;
   mapp<=66;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=17839;
 end   
19'd107703: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=89;
   mapp<=60;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10888;
 end   
19'd107704: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=94;
   mapp<=18;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=17453;
 end   
19'd107705: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=4;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd107706: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=19;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd107707: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd107708: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd107709: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd107710: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=65;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=35295;
 end   
19'd107711: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=24;
   mapp<=27;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=35917;
 end   
19'd107712: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=84;
   mapp<=88;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=37911;
 end   
19'd107713: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=25;
   mapp<=61;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=38235;
 end   
19'd107714: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=53;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd107715: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=92;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd107716: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd107717: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd107718: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd107719: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd107861: begin  
rid<=1;
end
19'd107862: begin  
end
19'd107863: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd107864: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd107865: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd107866: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd107867: begin  
rid<=0;
end
19'd108001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=56;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=21370;
 end   
19'd108002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=65;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=19176;
 end   
19'd108003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=36;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd108004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=69;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd108005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=24;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd108006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=86;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd108007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=72;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd108008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=2;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd108009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=52;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd108010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=71;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd108011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd108012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=93;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=52612;
 end   
19'd108013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=58;
   mapp<=25;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=49299;
 end   
19'd108014: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=40;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd108015: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=87;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd108016: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=88;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd108017: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=77;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd108018: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=59;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd108019: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=59;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd108020: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=30;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd108021: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=30;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd108022: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd108023: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd108165: begin  
rid<=1;
end
19'd108166: begin  
end
19'd108167: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd108168: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd108169: begin  
rid<=0;
end
19'd108301: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=60;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=15326;
 end   
19'd108302: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=94;
   mapp<=91;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12378;
 end   
19'd108303: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=28;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd108304: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=37;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd108305: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=53;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd108306: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=96;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=28166;
 end   
19'd108307: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=4;
   mapp<=39;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20062;
 end   
19'd108308: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=68;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd108309: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=96;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd108310: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=75;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd108311: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd108453: begin  
rid<=1;
end
19'd108454: begin  
end
19'd108455: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd108456: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd108457: begin  
rid<=0;
end
19'd108601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=1;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13994;
 end   
19'd108602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=7;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd108603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=95;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd108604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=52;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd108605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=35;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd108606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=60;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd108607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=52;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd108608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=63;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=36305;
 end   
19'd108609: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=12;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd108610: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=74;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd108611: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=49;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd108612: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=30;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd108613: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=28;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd108614: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=95;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd108615: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd108757: begin  
rid<=1;
end
19'd108758: begin  
end
19'd108759: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd108760: begin  
rid<=0;
end
19'd108901: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=45;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1215;
 end   
19'd108902: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10;
 end   
19'd108903: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=85;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2315;
 end   
19'd108904: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=90;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=2460;
 end   
19'd108905: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=72;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1984;
 end   
19'd108906: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=38;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=1076;
 end   
19'd108907: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=71;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=1977;
 end   
19'd108908: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=96;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=10143;
 end   
19'd108909: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=73;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=6799;
 end   
19'd108910: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=61;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=7988;
 end   
19'd108911: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=8;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=3204;
 end   
19'd108912: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=16;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=3472;
 end   
19'd108913: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=1076;
 end   
19'd108914: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=39;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=5604;
 end   
19'd108915: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd109057: begin  
rid<=1;
end
19'd109058: begin  
end
19'd109059: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd109060: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd109061: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd109062: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd109063: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd109064: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd109065: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd109066: begin  
rid<=0;
end
19'd109201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=72;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5184;
 end   
19'd109202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=78;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5626;
 end   
19'd109203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=89;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6428;
 end   
19'd109204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=78;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12438;
 end   
19'd109205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=58;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=10150;
 end   
19'd109206: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=99;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=14150;
 end   
19'd109207: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd109349: begin  
rid<=1;
end
19'd109350: begin  
end
19'd109351: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd109352: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd109353: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd109354: begin  
rid<=0;
end
19'd109501: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=26;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=30019;
 end   
19'd109502: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=94;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=31347;
 end   
19'd109503: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=45;
   mapp<=67;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=32337;
 end   
19'd109504: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=74;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd109505: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=48;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd109506: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=83;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd109507: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=44;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd109508: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=81;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd109509: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=75;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd109510: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd109511: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=91;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=49806;
 end   
19'd109512: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=89;
   mapp<=18;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=49506;
 end   
19'd109513: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=68;
   mapp<=98;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=49374;
 end   
19'd109514: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=60;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd109515: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=12;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd109516: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd109517: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=12;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd109518: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=34;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd109519: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=77;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd109520: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=75;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd109521: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd109663: begin  
rid<=1;
end
19'd109664: begin  
end
19'd109665: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd109666: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd109667: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd109668: begin  
rid<=0;
end
19'd109801: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=98;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4606;
 end   
19'd109802: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=90;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8830;
 end   
19'd109803: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=40;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3940;
 end   
19'd109804: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=5;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=520;
 end   
19'd109805: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=84;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=8272;
 end   
19'd109806: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=43;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=4264;
 end   
19'd109807: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=14;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=1432;
 end   
19'd109808: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=64;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=6342;
 end   
19'd109809: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=80;
 end   
19'd109810: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=60;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=9526;
 end   
19'd109811: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=75;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=13330;
 end   
19'd109812: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=8140;
 end   
19'd109813: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=23;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=1900;
 end   
19'd109814: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=98;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=14152;
 end   
19'd109815: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=51;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=7324;
 end   
19'd109816: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=64;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=5272;
 end   
19'd109817: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=77;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=10962;
 end   
19'd109818: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=23;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=1460;
 end   
19'd109819: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd109961: begin  
rid<=1;
end
19'd109962: begin  
end
19'd109963: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd109964: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd109965: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd109966: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd109967: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd109968: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd109969: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd109970: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd109971: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd109972: begin  
rid<=0;
end
19'd110101: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=13;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11812;
 end   
19'd110102: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=98;
   mapp<=70;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10925;
 end   
19'd110103: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=44;
   mapp<=19;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11518;
 end   
19'd110104: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=59;
   mapp<=55;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=15274;
 end   
19'd110105: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=97;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6807;
 end   
19'd110106: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=27;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=11963;
 end   
19'd110107: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=65;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=8848;
 end   
19'd110108: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd110109: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd110110: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd110111: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=87;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=18228;
 end   
19'd110112: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=31;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=16620;
 end   
19'd110113: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=64;
   mapp<=5;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=14068;
 end   
19'd110114: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=1;
   mapp<=10;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=17864;
 end   
19'd110115: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=28;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=11008;
 end   
19'd110116: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=13;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=18994;
 end   
19'd110117: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=20;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=15244;
 end   
19'd110118: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd110119: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd110120: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd110121: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd110263: begin  
rid<=1;
end
19'd110264: begin  
end
19'd110265: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd110266: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd110267: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd110268: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd110269: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd110270: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd110271: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd110272: begin  
rid<=0;
end
19'd110401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=94;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6823;
 end   
19'd110402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=27;
   mapp<=73;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9350;
 end   
19'd110403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=88;
   mapp<=53;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4244;
 end   
19'd110404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=54;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3782;
 end   
19'd110405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=2;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd110406: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=66;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd110407: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=37;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=11742;
 end   
19'd110408: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=33;
   mapp<=47;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=16560;
 end   
19'd110409: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=12;
   mapp<=71;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=9394;
 end   
19'd110410: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=62;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=9009;
 end   
19'd110411: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=20;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd110412: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=1;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd110413: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd110555: begin  
rid<=1;
end
19'd110556: begin  
end
19'd110557: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd110558: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd110559: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd110560: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd110561: begin  
rid<=0;
end
19'd110701: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=53;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=18953;
 end   
19'd110702: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=46;
   mapp<=17;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=16137;
 end   
19'd110703: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=13;
   mapp<=41;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=17338;
 end   
19'd110704: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=94;
   mapp<=63;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=20018;
 end   
19'd110705: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=7;
   mapp<=48;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=10776;
 end   
19'd110706: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=75;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd110707: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=66;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd110708: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=29;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd110709: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=82;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd110710: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=8;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd110711: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=2;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd110712: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=24;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=33223;
 end   
19'd110713: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=78;
   mapp<=71;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=30143;
 end   
19'd110714: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=1;
   mapp<=6;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=25370;
 end   
19'd110715: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=31;
   mapp<=98;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=36292;
 end   
19'd110716: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=40;
   mapp<=55;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=27884;
 end   
19'd110717: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=3;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd110718: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=25;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd110719: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=28;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd110720: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=59;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd110721: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd110722: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd110723: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd110865: begin  
rid<=1;
end
19'd110866: begin  
end
19'd110867: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd110868: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd110869: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd110870: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd110871: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd110872: begin  
rid<=0;
end
19'd111001: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2583;
 end   
19'd111002: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=41;
   mapp<=63;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4500;
 end   
19'd111003: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=14;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1567;
 end   
19'd111004: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=5;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3242;
 end   
19'd111005: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=44;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4605;
 end   
19'd111006: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=11;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=5743;
 end   
19'd111007: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=75;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd111008: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=58;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8037;
 end   
19'd111009: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=97;
   mapp<=6;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=13212;
 end   
19'd111010: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=94;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=9817;
 end   
19'd111011: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=59;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=8336;
 end   
19'd111012: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=23;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=6627;
 end   
19'd111013: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=15;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=7579;
 end   
19'd111014: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=96;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd111015: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd111157: begin  
rid<=1;
end
19'd111158: begin  
end
19'd111159: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd111160: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd111161: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd111162: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd111163: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd111164: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd111165: begin  
rid<=0;
end
19'd111301: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=5;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16195;
 end   
19'd111302: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=95;
   mapp<=76;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=17931;
 end   
19'd111303: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=87;
   mapp<=96;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=13809;
 end   
19'd111304: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=43;
   mapp<=6;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=10557;
 end   
19'd111305: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=41;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd111306: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=39;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd111307: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd111308: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=96;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=35785;
 end   
19'd111309: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=82;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=34224;
 end   
19'd111310: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=71;
   mapp<=72;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=29579;
 end   
19'd111311: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=85;
   mapp<=52;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=24597;
 end   
19'd111312: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=29;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd111313: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=84;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd111314: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=47;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd111315: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd111457: begin  
rid<=1;
end
19'd111458: begin  
end
19'd111459: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd111460: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd111461: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd111462: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd111463: begin  
rid<=0;
end
19'd111601: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=7;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1158;
 end   
19'd111602: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=31;
   mapp<=15;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=797;
 end   
19'd111603: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=22;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1476;
 end   
19'd111604: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=42;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=696;
 end   
19'd111605: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd111606: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=58;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5292;
 end   
19'd111607: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=25;
   mapp<=54;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=5704;
 end   
19'd111608: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=71;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=7844;
 end   
19'd111609: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=90;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6141;
 end   
19'd111610: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd111611: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd111753: begin  
rid<=1;
end
19'd111754: begin  
end
19'd111755: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd111756: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd111757: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd111758: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd111759: begin  
rid<=0;
end
19'd111901: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=84;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=17985;
 end   
19'd111902: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=26;
   mapp<=55;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=22110;
 end   
19'd111903: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=86;
   mapp<=5;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10577;
 end   
19'd111904: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=11;
   mapp<=89;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=20025;
 end   
19'd111905: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=22;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd111906: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=69;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd111907: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=58;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd111908: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=11;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd111909: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd111910: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd111911: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd111912: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=47;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=33850;
 end   
19'd111913: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=19;
   mapp<=4;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=28842;
 end   
19'd111914: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=91;
   mapp<=85;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=25530;
 end   
19'd111915: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=48;
   mapp<=3;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=27538;
 end   
19'd111916: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=60;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd111917: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=5;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd111918: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=25;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd111919: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=90;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd111920: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd111921: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd111922: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd111923: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd112065: begin  
rid<=1;
end
19'd112066: begin  
end
19'd112067: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd112068: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd112069: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd112070: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd112071: begin  
rid<=0;
end
19'd112201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=11;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10734;
 end   
19'd112202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=84;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd112203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=47;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd112204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=0;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=15099;
 end   
19'd112205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=61;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd112206: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=17;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd112207: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd112349: begin  
rid<=1;
end
19'd112350: begin  
end
19'd112351: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd112352: begin  
rid<=0;
end
19'd112501: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=85;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4988;
 end   
19'd112502: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=89;
   mapp<=23;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5488;
 end   
19'd112503: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=7;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd112504: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=44;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd112505: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=35;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd112506: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=64;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd112507: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=12;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd112508: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=27;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd112509: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=15;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=19955;
 end   
19'd112510: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=41;
   mapp<=55;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20801;
 end   
19'd112511: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=56;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd112512: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=9;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd112513: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=19;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd112514: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=27;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd112515: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=62;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd112516: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=48;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd112517: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd112659: begin  
rid<=1;
end
19'd112660: begin  
end
19'd112661: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd112662: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd112663: begin  
rid<=0;
end
19'd112801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=6;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4878;
 end   
19'd112802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=91;
   mapp<=51;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5053;
 end   
19'd112803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=1;
   mapp<=51;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9160;
 end   
19'd112804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=96;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=9603;
 end   
19'd112805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=98;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=7855;
 end   
19'd112806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd112807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd112808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=41;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=11651;
 end   
19'd112809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=55;
   mapp<=81;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=13594;
 end   
19'd112810: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=35;
   mapp<=51;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=18056;
 end   
19'd112811: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=69;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=19857;
 end   
19'd112812: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=86;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=17086;
 end   
19'd112813: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd112814: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd112815: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd112957: begin  
rid<=1;
end
19'd112958: begin  
end
19'd112959: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd112960: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd112961: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd112962: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd112963: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd112964: begin  
rid<=0;
end
19'd113101: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=56;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=23400;
 end   
19'd113102: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=93;
   mapp<=80;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=20605;
 end   
19'd113103: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=73;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd113104: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=71;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd113105: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=31;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd113106: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd113107: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=37064;
 end   
19'd113108: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=66;
   mapp<=53;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=31559;
 end   
19'd113109: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=92;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd113110: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=46;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd113111: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=64;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd113112: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd113113: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd113255: begin  
rid<=1;
end
19'd113256: begin  
end
19'd113257: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd113258: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd113259: begin  
rid<=0;
end
19'd113401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=65;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3425;
 end   
19'd113402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=5;
   mapp<=9;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=760;
 end   
19'd113403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=33;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2275;
 end   
19'd113404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=22;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1870;
 end   
19'd113405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=82;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5815;
 end   
19'd113406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=89;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6045;
 end   
19'd113407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=42;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=2810;
 end   
19'd113408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=4;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=675;
 end   
19'd113409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=69;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=4765;
 end   
19'd113410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=40;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=2870;
 end   
19'd113411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd113412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=13;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=10493;
 end   
19'd113413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=96;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=4192;
 end   
19'd113414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=26;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=7893;
 end   
19'd113415: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=55;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=4985;
 end   
19'd113416: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=25;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=7100;
 end   
19'd113417: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=10;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=11551;
 end   
19'd113418: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=56;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=11986;
 end   
19'd113419: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=88;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=6235;
 end   
19'd113420: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=46;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=11891;
 end   
19'd113421: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=68;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=5098;
 end   
19'd113422: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd113423: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd113565: begin  
rid<=1;
end
19'd113566: begin  
end
19'd113567: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd113568: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd113569: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd113570: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd113571: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd113572: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd113573: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd113574: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd113575: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd113576: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd113577: begin  
rid<=0;
end
19'd113701: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=56;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12352;
 end   
19'd113702: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=88;
   mapp<=81;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9888;
 end   
19'd113703: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=16;
   mapp<=29;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7300;
 end   
19'd113704: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=38;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=11633;
 end   
19'd113705: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=98;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=12456;
 end   
19'd113706: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=15;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=9982;
 end   
19'd113707: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=99;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd113708: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=22;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd113709: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=43;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=15671;
 end   
19'd113710: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=16;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=14089;
 end   
19'd113711: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=28;
   mapp<=29;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=14982;
 end   
19'd113712: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=61;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=20462;
 end   
19'd113713: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=90;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=18247;
 end   
19'd113714: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=24;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=14925;
 end   
19'd113715: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=41;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd113716: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=47;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd113717: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd113859: begin  
rid<=1;
end
19'd113860: begin  
end
19'd113861: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd113862: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd113863: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd113864: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd113865: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd113866: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd113867: begin  
rid<=0;
end
19'd114001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=49;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=19923;
 end   
19'd114002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=90;
   mapp<=82;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=21090;
 end   
19'd114003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=91;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd114004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=68;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd114005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=45;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd114006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=17;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd114007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=25;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=32940;
 end   
19'd114008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=2;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=39118;
 end   
19'd114009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=82;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd114010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=95;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd114011: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=28;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd114012: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=55;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd114013: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd114155: begin  
rid<=1;
end
19'd114156: begin  
end
19'd114157: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd114158: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd114159: begin  
rid<=0;
end
19'd114301: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=65;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=21228;
 end   
19'd114302: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=97;
   mapp<=13;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=17807;
 end   
19'd114303: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=68;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd114304: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=16;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd114305: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=18;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd114306: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=44;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd114307: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=4;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd114308: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=63;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd114309: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=79;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd114310: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=15;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd114311: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=36;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=36247;
 end   
19'd114312: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=58;
   mapp<=43;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=36038;
 end   
19'd114313: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd114314: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=22;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd114315: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=74;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd114316: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=35;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd114317: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=28;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd114318: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=14;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd114319: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=58;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd114320: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=99;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd114321: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd114463: begin  
rid<=1;
end
19'd114464: begin  
end
19'd114465: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd114466: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd114467: begin  
rid<=0;
end
19'd114601: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=18;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=458;
 end   
19'd114602: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=2;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=908;
 end   
19'd114603: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=89;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1694;
 end   
19'd114604: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=36;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=764;
 end   
19'd114605: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=43;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1000;
 end   
19'd114606: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=93;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=1816;
 end   
19'd114607: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=46;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=930;
 end   
19'd114608: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=21;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=504;
 end   
19'd114609: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=28;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=772;
 end   
19'd114610: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd114611: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=66;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8480;
 end   
19'd114612: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=54;
   mapp<=96;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8702;
 end   
19'd114613: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=27;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=4394;
 end   
19'd114614: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=17;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6476;
 end   
19'd114615: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=85;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=6772;
 end   
19'd114616: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=3;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=5902;
 end   
19'd114617: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=72;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=9786;
 end   
19'd114618: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=76;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=10110;
 end   
19'd114619: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=85;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=6976;
 end   
19'd114620: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd114621: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd114763: begin  
rid<=1;
end
19'd114764: begin  
end
19'd114765: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd114766: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd114767: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd114768: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd114769: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd114770: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd114771: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd114772: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd114773: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd114774: begin  
rid<=0;
end
19'd114901: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=9;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5287;
 end   
19'd114902: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=34;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6884;
 end   
19'd114903: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=98;
   mapp<=50;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9390;
 end   
19'd114904: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=0;
   mapp<=66;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6440;
 end   
19'd114905: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=82;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=13954;
 end   
19'd114906: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=16;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=8886;
 end   
19'd114907: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=85;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=7949;
 end   
19'd114908: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=93;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd114909: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=53;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd114910: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=24;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd114911: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=43;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7787;
 end   
19'd114912: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=3;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=9952;
 end   
19'd114913: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=23;
   mapp<=11;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=17269;
 end   
19'd114914: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=16;
   mapp<=75;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=9040;
 end   
19'd114915: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=23;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=19450;
 end   
19'd114916: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=85;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=12222;
 end   
19'd114917: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=3;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=15075;
 end   
19'd114918: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd114919: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=17;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd114920: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=84;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd114921: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd115063: begin  
rid<=1;
end
19'd115064: begin  
end
19'd115065: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd115066: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd115067: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd115068: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd115069: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd115070: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd115071: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd115072: begin  
rid<=0;
end
19'd115201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=65;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4290;
 end   
19'd115202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=4;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=270;
 end   
19'd115203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=84;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5480;
 end   
19'd115204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=81;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5295;
 end   
19'd115205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=15;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5370;
 end   
19'd115206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=30;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=720;
 end   
19'd115207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=60;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=6380;
 end   
19'd115208: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=87;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6600;
 end   
19'd115209: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd115351: begin  
rid<=1;
end
19'd115352: begin  
end
19'd115353: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd115354: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd115355: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd115356: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd115357: begin  
rid<=0;
end
19'd115501: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=67;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1407;
 end   
19'd115502: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=42;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2824;
 end   
19'd115503: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=65;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4375;
 end   
19'd115504: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=49;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3313;
 end   
19'd115505: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=58;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3926;
 end   
19'd115506: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=48;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=3266;
 end   
19'd115507: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=66;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=4482;
 end   
19'd115508: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=70;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=4760;
 end   
19'd115509: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=96;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=6512;
 end   
19'd115510: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=93;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=6321;
 end   
19'd115511: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=3;
   pp<=100;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[10]<=301;
 end   
19'd115512: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=72;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7383;
 end   
19'd115513: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=60;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=7144;
 end   
19'd115514: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=14;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=5383;
 end   
19'd115515: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=44;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6481;
 end   
19'd115516: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=15;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=5006;
 end   
19'd115517: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=14;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=4274;
 end   
19'd115518: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=24;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=6210;
 end   
19'd115519: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=61;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=9152;
 end   
19'd115520: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=25;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=8312;
 end   
19'd115521: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=6321;
 end   
19'd115522: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=67;
   pp<=100;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[10]<=5125;
 end   
19'd115523: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd115665: begin  
rid<=1;
end
19'd115666: begin  
end
19'd115667: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd115668: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd115669: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd115670: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd115671: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd115672: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd115673: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd115674: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd115675: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd115676: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd115677: begin  
check0<=expctdoutput[10]-outcheck0;
end
19'd115678: begin  
rid<=0;
end
19'd115801: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=79;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1422;
 end   
19'd115802: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=13;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1037;
 end   
19'd115803: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=58;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4602;
 end   
19'd115804: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=24;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=3078;
 end   
19'd115805: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=86;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=3101;
 end   
19'd115806: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=75;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=6402;
 end   
19'd115807: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd115949: begin  
rid<=1;
end
19'd115950: begin  
end
19'd115951: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd115952: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd115953: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd115954: begin  
rid<=0;
end
19'd116101: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=82;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1394;
 end   
19'd116102: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=71;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1217;
 end   
19'd116103: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=40;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=700;
 end   
19'd116104: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=1;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=47;
 end   
19'd116105: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=35;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=635;
 end   
19'd116106: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=25;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=475;
 end   
19'd116107: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=73;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=1301;
 end   
19'd116108: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=6;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=1676;
 end   
19'd116109: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=88;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=5353;
 end   
19'd116110: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=17;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=1499;
 end   
19'd116111: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=43;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=2068;
 end   
19'd116112: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=38;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=2421;
 end   
19'd116113: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=84;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=4423;
 end   
19'd116114: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=57;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=3980;
 end   
19'd116115: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd116257: begin  
rid<=1;
end
19'd116258: begin  
end
19'd116259: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd116260: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd116261: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd116262: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd116263: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd116264: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd116265: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd116266: begin  
rid<=0;
end
19'd116401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=91;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=25622;
 end   
19'd116402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=99;
   mapp<=31;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=35236;
 end   
19'd116403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=91;
   mapp<=53;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=33870;
 end   
19'd116404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=40;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd116405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=90;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd116406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=6;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd116407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=13;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd116408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=98;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd116409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=23;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd116410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd116411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd116412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=98;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=54021;
 end   
19'd116413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=46;
   mapp<=62;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=58489;
 end   
19'd116414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=87;
   mapp<=25;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=53243;
 end   
19'd116415: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=78;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd116416: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=12;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd116417: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=18;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd116418: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=82;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd116419: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=84;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd116420: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=14;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd116421: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd116422: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd116423: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd116565: begin  
rid<=1;
end
19'd116566: begin  
end
19'd116567: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd116568: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd116569: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd116570: begin  
rid<=0;
end
19'd116701: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=92;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9312;
 end   
19'd116702: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=66;
   mapp<=27;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5913;
 end   
19'd116703: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=24;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd116704: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=44;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd116705: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=55;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd116706: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=2;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd116707: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=35;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=25215;
 end   
19'd116708: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=68;
   mapp<=88;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=17478;
 end   
19'd116709: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=99;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd116710: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=10;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd116711: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=13;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd116712: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=8;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd116713: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd116855: begin  
rid<=1;
end
19'd116856: begin  
end
19'd116857: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd116858: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd116859: begin  
rid<=0;
end
19'd117001: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=92;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12937;
 end   
19'd117002: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=84;
   mapp<=54;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10606;
 end   
19'd117003: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=81;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd117004: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=48;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd117005: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=40;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd117006: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=24;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd117007: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=1;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd117008: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd117009: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=78;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=32728;
 end   
19'd117010: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=14;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=23297;
 end   
19'd117011: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=7;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd117012: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=73;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd117013: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=99;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd117014: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=66;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd117015: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=68;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd117016: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd117017: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd117159: begin  
rid<=1;
end
19'd117160: begin  
end
19'd117161: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd117162: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd117163: begin  
rid<=0;
end
19'd117301: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=88;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=28176;
 end   
19'd117302: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=72;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd117303: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=38;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd117304: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=13;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd117305: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=33;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd117306: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=48;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd117307: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=31;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd117308: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=50;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd117309: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=96;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd117310: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=59;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd117311: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=9;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd117312: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=39;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=50772;
 end   
19'd117313: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=7;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd117314: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=29;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd117315: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=13;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd117316: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=54;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd117317: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=85;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd117318: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=50;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd117319: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=93;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd117320: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=49;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd117321: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=94;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd117322: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=2;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd117323: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd117465: begin  
rid<=1;
end
19'd117466: begin  
end
19'd117467: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd117468: begin  
rid<=0;
end
19'd117601: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=96;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5616;
 end   
19'd117602: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=42;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7216;
 end   
19'd117603: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd117604: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=19;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8034;
 end   
19'd117605: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=21;
   mapp<=50;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8334;
 end   
19'd117606: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd117607: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd117749: begin  
rid<=1;
end
19'd117750: begin  
end
19'd117751: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd117752: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd117753: begin  
rid<=0;
end
19'd117901: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=58;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4609;
 end   
19'd117902: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=75;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3600;
 end   
19'd117903: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd117904: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=52;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14450;
 end   
19'd117905: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=83;
   mapp<=91;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=11154;
 end   
19'd117906: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd117907: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd118049: begin  
rid<=1;
end
19'd118050: begin  
end
19'd118051: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd118052: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd118053: begin  
rid<=0;
end
19'd118201: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=28;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3936;
 end   
19'd118202: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=51;
   mapp<=31;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4712;
 end   
19'd118203: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=61;
   mapp<=1;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6366;
 end   
19'd118204: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=10;
   mapp<=53;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6865;
 end   
19'd118205: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd118206: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd118207: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd118208: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=26;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16324;
 end   
19'd118209: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=69;
   mapp<=53;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=16780;
 end   
19'd118210: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=34;
   mapp<=27;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=19717;
 end   
19'd118211: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=63;
   mapp<=91;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=17845;
 end   
19'd118212: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd118213: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd118214: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd118215: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd118357: begin  
rid<=1;
end
19'd118358: begin  
end
19'd118359: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd118360: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd118361: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd118362: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd118363: begin  
rid<=0;
end
19'd118501: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=11;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1962;
 end   
19'd118502: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=25;
   mapp<=49;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=974;
 end   
19'd118503: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=17;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1832;
 end   
19'd118504: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd118505: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=15;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8220;
 end   
19'd118506: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=99;
   mapp<=62;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=6854;
 end   
19'd118507: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=50;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=4958;
 end   
19'd118508: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd118509: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd118651: begin  
rid<=1;
end
19'd118652: begin  
end
19'd118653: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd118654: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd118655: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd118656: begin  
rid<=0;
end
19'd118801: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=7;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9496;
 end   
19'd118802: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=35;
   mapp<=21;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11747;
 end   
19'd118803: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=66;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd118804: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=92;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd118805: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd118806: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=44;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=19990;
 end   
19'd118807: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=70;
   mapp<=49;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20661;
 end   
19'd118808: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=59;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd118809: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=33;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd118810: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=0;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd118811: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd118953: begin  
rid<=1;
end
19'd118954: begin  
end
19'd118955: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd118956: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd118957: begin  
rid<=0;
end
19'd119101: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=74;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=28754;
 end   
19'd119102: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=89;
   mapp<=22;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=25605;
 end   
19'd119103: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=59;
   mapp<=5;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=25941;
 end   
19'd119104: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=64;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd119105: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=79;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd119106: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=72;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd119107: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=69;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd119108: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=8;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd119109: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=17;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd119110: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd119111: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd119112: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=24;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=57417;
 end   
19'd119113: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=26;
   mapp<=22;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=54992;
 end   
19'd119114: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=63;
   mapp<=18;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=52359;
 end   
19'd119115: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=91;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd119116: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=92;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd119117: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=92;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd119118: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=54;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd119119: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=30;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd119120: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=49;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd119121: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd119122: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd119123: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd119265: begin  
rid<=1;
end
19'd119266: begin  
end
19'd119267: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd119268: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd119269: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd119270: begin  
rid<=0;
end
19'd119401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=71;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12450;
 end   
19'd119402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=37;
   mapp<=91;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12547;
 end   
19'd119403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=40;
   mapp<=62;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=15096;
 end   
19'd119404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=88;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=17034;
 end   
19'd119405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=54;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=14949;
 end   
19'd119406: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=63;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd119407: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=67;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd119408: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=13;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14899;
 end   
19'd119409: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=6;
   mapp<=61;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18898;
 end   
19'd119410: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=85;
   mapp<=19;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=21282;
 end   
19'd119411: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=50;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=19838;
 end   
19'd119412: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=4;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=18901;
 end   
19'd119413: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=40;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd119414: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=72;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd119415: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd119557: begin  
rid<=1;
end
19'd119558: begin  
end
19'd119559: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd119560: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd119561: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd119562: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd119563: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd119564: begin  
rid<=0;
end
19'd119701: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=96;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4320;
 end   
19'd119702: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=6;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=586;
 end   
19'd119703: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=26;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2516;
 end   
19'd119704: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=57;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5502;
 end   
19'd119705: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=93;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8598;
 end   
19'd119706: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=80;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8026;
 end   
19'd119707: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=96;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=11444;
 end   
19'd119708: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=84;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=13314;
 end   
19'd119709: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd119851: begin  
rid<=1;
end
19'd119852: begin  
end
19'd119853: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd119854: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd119855: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd119856: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd119857: begin  
rid<=0;
end
19'd120001: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=56;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6306;
 end   
19'd120002: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=79;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd120003: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=29;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=13682;
 end   
19'd120004: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=56;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd120005: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd120147: begin  
rid<=1;
end
19'd120148: begin  
end
19'd120149: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd120150: begin  
rid<=0;
end
19'd120301: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=79;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2844;
 end   
19'd120302: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=94;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3394;
 end   
19'd120303: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=43;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1568;
 end   
19'd120304: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=6;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=246;
 end   
19'd120305: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=32;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1192;
 end   
19'd120306: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=79;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=2894;
 end   
19'd120307: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=90;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=3300;
 end   
19'd120308: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=81;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5679;
 end   
19'd120309: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=16;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=3954;
 end   
19'd120310: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=77;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=4263;
 end   
19'd120311: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=73;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=2801;
 end   
19'd120312: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=17;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=1787;
 end   
19'd120313: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=78;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=5624;
 end   
19'd120314: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=3;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=3405;
 end   
19'd120315: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd120457: begin  
rid<=1;
end
19'd120458: begin  
end
19'd120459: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd120460: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd120461: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd120462: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd120463: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd120464: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd120465: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd120466: begin  
rid<=0;
end
19'd120601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=9;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6398;
 end   
19'd120602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=35;
   mapp<=75;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7490;
 end   
19'd120603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=21;
   mapp<=32;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8164;
 end   
19'd120604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=37;
   mapp<=40;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=9709;
 end   
19'd120605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=43;
   mapp<=31;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=10478;
 end   
19'd120606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd120607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd120608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd120609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd120610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=7;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14518;
 end   
19'd120611: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=52;
   mapp<=6;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20882;
 end   
19'd120612: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=26;
   mapp<=96;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=18827;
 end   
19'd120613: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=31;
   mapp<=86;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=15566;
 end   
19'd120614: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=69;
   mapp<=35;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=15896;
 end   
19'd120615: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd120616: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd120617: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd120618: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd120619: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd120761: begin  
rid<=1;
end
19'd120762: begin  
end
19'd120763: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd120764: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd120765: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd120766: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd120767: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd120768: begin  
rid<=0;
end
19'd120901: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=30;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13986;
 end   
19'd120902: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=61;
   mapp<=7;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11762;
 end   
19'd120903: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=47;
   mapp<=46;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=14407;
 end   
19'd120904: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=70;
   mapp<=78;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=11313;
 end   
19'd120905: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=26;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd120906: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=87;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd120907: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=14;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd120908: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=86;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd120909: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=5;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd120910: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=20;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=20652;
 end   
19'd120911: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=16;
   mapp<=65;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=21690;
 end   
19'd120912: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=38;
   mapp<=21;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=23761;
 end   
19'd120913: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=31;
   mapp<=44;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=21009;
 end   
19'd120914: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=88;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd120915: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=44;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd120916: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=39;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd120917: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=35;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd120918: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=1;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd120919: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd121061: begin  
rid<=1;
end
19'd121062: begin  
end
19'd121063: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd121064: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd121065: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd121066: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd121067: begin  
rid<=0;
end
19'd121201: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=86;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8495;
 end   
19'd121202: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=28;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6588;
 end   
19'd121203: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=9;
   mapp<=34;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6617;
 end   
19'd121204: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=63;
   mapp<=41;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6690;
 end   
19'd121205: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=0;
   mapp<=65;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6622;
 end   
19'd121206: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=5;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd121207: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=30;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd121208: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=31;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd121209: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=10;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd121210: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=5;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd121211: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=97;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd121212: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=11;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=22691;
 end   
19'd121213: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=60;
   mapp<=16;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=21381;
 end   
19'd121214: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=35;
   mapp<=96;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=17761;
 end   
19'd121215: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=90;
   mapp<=89;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=21626;
 end   
19'd121216: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=20;
   mapp<=33;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=21473;
 end   
19'd121217: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=46;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd121218: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=60;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd121219: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=45;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd121220: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=90;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd121221: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=45;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd121222: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd121223: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd121365: begin  
rid<=1;
end
19'd121366: begin  
end
19'd121367: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd121368: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd121369: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd121370: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd121371: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd121372: begin  
rid<=0;
end
19'd121501: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=56;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1102;
 end   
19'd121502: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=1;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4377;
 end   
19'd121503: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=79;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd121504: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd121505: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=46;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8112;
 end   
19'd121506: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=43;
   mapp<=54;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8161;
 end   
19'd121507: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=14;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd121508: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd121509: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd121651: begin  
rid<=1;
end
19'd121652: begin  
end
19'd121653: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd121654: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd121655: begin  
rid<=0;
end
19'd121801: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=60;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=15702;
 end   
19'd121802: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=30;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9484;
 end   
19'd121803: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=11;
   mapp<=69;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=13753;
 end   
19'd121804: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=9;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd121805: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=68;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd121806: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=30;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd121807: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=38;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd121808: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=32;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd121809: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=1;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd121810: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=2;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd121811: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=91;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd121812: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=49;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=32410;
 end   
19'd121813: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=12;
   mapp<=4;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=24867;
 end   
19'd121814: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=46;
   mapp<=79;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=31954;
 end   
19'd121815: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=18;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd121816: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=38;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd121817: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=89;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd121818: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=90;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd121819: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=33;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd121820: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=72;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd121821: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd121822: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=53;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd121823: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd121965: begin  
rid<=1;
end
19'd121966: begin  
end
19'd121967: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd121968: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd121969: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd121970: begin  
rid<=0;
end
19'd122101: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=68;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4450;
 end   
19'd122102: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=37;
   mapp<=70;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8259;
 end   
19'd122103: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=24;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd122104: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd122105: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=58;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16586;
 end   
19'd122106: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=86;
   mapp<=88;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20959;
 end   
19'd122107: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=20;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd122108: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd122109: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd122251: begin  
rid<=1;
end
19'd122252: begin  
end
19'd122253: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd122254: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd122255: begin  
rid<=0;
end
19'd122401: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=89;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13076;
 end   
19'd122402: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=83;
   mapp<=9;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11073;
 end   
19'd122403: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=21;
   mapp<=91;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=19615;
 end   
19'd122404: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=87;
   mapp<=42;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=8121;
 end   
19'd122405: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd122406: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd122407: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd122408: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=6;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=15656;
 end   
19'd122409: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=19;
   mapp<=24;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12665;
 end   
19'd122410: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=43;
   mapp<=38;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=22885;
 end   
19'd122411: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=2;
   mapp<=14;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=11902;
 end   
19'd122412: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd122413: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd122414: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd122415: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd122557: begin  
rid<=1;
end
19'd122558: begin  
end
19'd122559: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd122560: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd122561: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd122562: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd122563: begin  
rid<=0;
end
19'd122701: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=48;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6867;
 end   
19'd122702: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=15;
   mapp<=7;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4433;
 end   
19'd122703: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=79;
   mapp<=18;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10543;
 end   
19'd122704: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=21;
   mapp<=44;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7044;
 end   
19'd122705: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=48;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=9679;
 end   
19'd122706: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=51;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=10177;
 end   
19'd122707: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=87;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=12563;
 end   
19'd122708: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=75;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=12219;
 end   
19'd122709: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=79;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd122710: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=58;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd122711: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=83;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd122712: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=25;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=18462;
 end   
19'd122713: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=95;
   mapp<=87;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=22083;
 end   
19'd122714: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=60;
   mapp<=7;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=21569;
 end   
19'd122715: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=20;
   mapp<=88;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=21191;
 end   
19'd122716: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=90;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=24792;
 end   
19'd122717: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=67;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=24845;
 end   
19'd122718: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=56;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=24389;
 end   
19'd122719: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=54;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=26217;
 end   
19'd122720: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=72;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd122721: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=46;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd122722: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=56;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd122723: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd122865: begin  
rid<=1;
end
19'd122866: begin  
end
19'd122867: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd122868: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd122869: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd122870: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd122871: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd122872: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd122873: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd122874: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd122875: begin  
rid<=0;
end
19'd123001: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=9;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=861;
 end   
19'd123002: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=8;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd123003: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=71;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14016;
 end   
19'd123004: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=80;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd123005: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd123147: begin  
rid<=1;
end
19'd123148: begin  
end
19'd123149: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd123150: begin  
rid<=0;
end
19'd123301: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=57;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7869;
 end   
19'd123302: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=21;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7466;
 end   
19'd123303: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=56;
   mapp<=93;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11092;
 end   
19'd123304: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=3;
   mapp<=94;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=11161;
 end   
19'd123305: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=66;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=12114;
 end   
19'd123306: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=28;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd123307: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd123308: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd123309: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=20;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=10947;
 end   
19'd123310: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=2;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=11318;
 end   
19'd123311: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=2;
   mapp<=72;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=13761;
 end   
19'd123312: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=48;
   mapp<=33;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=17392;
 end   
19'd123313: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=6;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=17675;
 end   
19'd123314: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=13;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd123315: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=61;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd123316: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=10;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd123317: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd123459: begin  
rid<=1;
end
19'd123460: begin  
end
19'd123461: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd123462: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd123463: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd123464: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd123465: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd123466: begin  
rid<=0;
end
19'd123601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=88;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12734;
 end   
19'd123602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=74;
   mapp<=71;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=13066;
 end   
19'd123603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=92;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9004;
 end   
19'd123604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=12;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3898;
 end   
19'd123605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=38;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=9970;
 end   
19'd123606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=89;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7956;
 end   
19'd123607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=1;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=5254;
 end   
19'd123608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=69;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=6808;
 end   
19'd123609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd123610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=20;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14817;
 end   
19'd123611: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=9;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=14748;
 end   
19'd123612: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=38;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=10268;
 end   
19'd123613: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=56;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=5900;
 end   
19'd123614: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=98;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=12182;
 end   
19'd123615: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=28;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=8993;
 end   
19'd123616: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=53;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=6395;
 end   
19'd123617: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=9;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=7564;
 end   
19'd123618: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd123619: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd123761: begin  
rid<=1;
end
19'd123762: begin  
end
19'd123763: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd123764: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd123765: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd123766: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd123767: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd123768: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd123769: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd123770: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd123771: begin  
rid<=0;
end
19'd123901: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=39;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13732;
 end   
19'd123902: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=40;
   mapp<=18;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12279;
 end   
19'd123903: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=19;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd123904: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=80;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd123905: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=93;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd123906: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=57;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd123907: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=92;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd123908: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=26;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd123909: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd123910: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=89;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=43334;
 end   
19'd123911: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=80;
   mapp<=39;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=39322;
 end   
19'd123912: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=65;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd123913: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=83;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd123914: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=94;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd123915: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=63;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd123916: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=13;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd123917: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=25;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd123918: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=61;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd123919: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd124061: begin  
rid<=1;
end
19'd124062: begin  
end
19'd124063: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd124064: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd124065: begin  
rid<=0;
end
19'd124201: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=92;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=17793;
 end   
19'd124202: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=50;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=20095;
 end   
19'd124203: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=85;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd124204: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=20;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd124205: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=31;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd124206: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=16;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd124207: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=86;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd124208: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd124209: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=34;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=40494;
 end   
19'd124210: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=23;
   mapp<=91;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=44505;
 end   
19'd124211: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=72;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd124212: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=48;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd124213: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=23;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd124214: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=91;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd124215: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=66;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd124216: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd124217: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd124359: begin  
rid<=1;
end
19'd124360: begin  
end
19'd124361: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd124362: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd124363: begin  
rid<=0;
end
19'd124501: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=61;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2501;
 end   
19'd124502: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=43;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1773;
 end   
19'd124503: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=45;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1865;
 end   
19'd124504: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=96;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3966;
 end   
19'd124505: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=29;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1229;
 end   
19'd124506: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=73;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=3043;
 end   
19'd124507: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=60;
 end   
19'd124508: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=50;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=2120;
 end   
19'd124509: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=3;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=203;
 end   
19'd124510: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=28;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=1238;
 end   
19'd124511: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=41;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=3772;
 end   
19'd124512: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=23;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=2486;
 end   
19'd124513: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=42;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=3167;
 end   
19'd124514: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=10;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=4276;
 end   
19'd124515: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=88;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=3957;
 end   
19'd124516: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=13;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=3446;
 end   
19'd124517: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=88;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=2788;
 end   
19'd124518: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=79;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=4569;
 end   
19'd124519: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=73;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=2466;
 end   
19'd124520: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=20;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=1858;
 end   
19'd124521: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd124663: begin  
rid<=1;
end
19'd124664: begin  
end
19'd124665: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd124666: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd124667: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd124668: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd124669: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd124670: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd124671: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd124672: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd124673: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd124674: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd124675: begin  
rid<=0;
end
19'd124801: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=31;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=434;
 end   
19'd124802: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10;
 end   
19'd124803: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=97;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1378;
 end   
19'd124804: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=8;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=522;
 end   
19'd124805: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=17;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=197;
 end   
19'd124806: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=2;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=1400;
 end   
19'd124807: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd124949: begin  
rid<=1;
end
19'd124950: begin  
end
19'd124951: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd124952: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd124953: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd124954: begin  
rid<=0;
end
19'd125101: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=96;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13704;
 end   
19'd125102: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=84;
   mapp<=29;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=13618;
 end   
19'd125103: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=76;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd125104: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd125105: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=3;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14908;
 end   
19'd125106: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=64;
   mapp<=13;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=22494;
 end   
19'd125107: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=95;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd125108: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd125109: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd125251: begin  
rid<=1;
end
19'd125252: begin  
end
19'd125253: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd125254: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd125255: begin  
rid<=0;
end
19'd125401: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=60;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13418;
 end   
19'd125402: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=89;
   mapp<=45;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=13355;
 end   
19'd125403: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=70;
   mapp<=64;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=13595;
 end   
19'd125404: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=49;
   mapp<=22;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=13487;
 end   
19'd125405: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=97;
   mapp<=15;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=11010;
 end   
19'd125406: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=91;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd125407: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=24;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd125408: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=52;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd125409: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=21;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd125410: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=96;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=24877;
 end   
19'd125411: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=48;
   mapp<=13;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=26034;
 end   
19'd125412: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=64;
   mapp<=35;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=26830;
 end   
19'd125413: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=58;
   mapp<=16;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=21104;
 end   
19'd125414: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=43;
   mapp<=89;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=19899;
 end   
19'd125415: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=81;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd125416: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=80;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd125417: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=7;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd125418: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=36;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd125419: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd125561: begin  
rid<=1;
end
19'd125562: begin  
end
19'd125563: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd125564: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd125565: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd125566: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd125567: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd125568: begin  
rid<=0;
end
19'd125701: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=31;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=18640;
 end   
19'd125702: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=61;
   mapp<=66;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=19937;
 end   
19'd125703: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd125704: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=93;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd125705: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=41;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd125706: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=49;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd125707: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=44;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd125708: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=10;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=28854;
 end   
19'd125709: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=42;
   mapp<=82;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=29256;
 end   
19'd125710: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=19;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd125711: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=13;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd125712: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=80;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd125713: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=8;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd125714: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=6;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd125715: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd125857: begin  
rid<=1;
end
19'd125858: begin  
end
19'd125859: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd125860: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd125861: begin  
rid<=0;
end
19'd126001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=56;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7207;
 end   
19'd126002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=35;
   mapp<=96;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15531;
 end   
19'd126003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=11;
   mapp<=71;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10857;
 end   
19'd126004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=87;
   mapp<=0;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=17101;
 end   
19'd126005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=2;
   mapp<=77;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=10842;
 end   
19'd126006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=84;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=14983;
 end   
19'd126007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=23;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=16230;
 end   
19'd126008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=83;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd126009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=13;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd126010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=32;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd126011: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=79;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd126012: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=7;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=13081;
 end   
19'd126013: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=9;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=22145;
 end   
19'd126014: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=15;
   mapp<=16;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=17474;
 end   
19'd126015: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=65;
   mapp<=58;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=27063;
 end   
19'd126016: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=30;
   mapp<=43;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=20421;
 end   
19'd126017: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=72;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=29609;
 end   
19'd126018: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=17;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=25547;
 end   
19'd126019: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=58;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd126020: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=81;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd126021: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=72;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd126022: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=57;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd126023: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd126165: begin  
rid<=1;
end
19'd126166: begin  
end
19'd126167: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd126168: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd126169: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd126170: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd126171: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd126172: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd126173: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd126174: begin  
rid<=0;
end
19'd126301: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=98;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=27154;
 end   
19'd126302: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=82;
   mapp<=11;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=31003;
 end   
19'd126303: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=52;
   mapp<=57;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=32040;
 end   
19'd126304: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=77;
   mapp<=93;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=35031;
 end   
19'd126305: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=57;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd126306: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=85;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd126307: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=93;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd126308: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd126309: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd126310: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd126311: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=77;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=45907;
 end   
19'd126312: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=27;
   mapp<=28;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=46838;
 end   
19'd126313: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=5;
   mapp<=94;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=47204;
 end   
19'd126314: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=91;
   mapp<=91;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=56193;
 end   
19'd126315: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=91;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd126316: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=83;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd126317: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=81;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd126318: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd126319: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd126320: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd126321: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd126463: begin  
rid<=1;
end
19'd126464: begin  
end
19'd126465: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd126466: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd126467: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd126468: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd126469: begin  
rid<=0;
end
19'd126601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=37;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14977;
 end   
19'd126602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=88;
   mapp<=18;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=16624;
 end   
19'd126603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=55;
   mapp<=14;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=15273;
 end   
19'd126604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=77;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd126605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=51;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd126606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=68;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd126607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=84;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd126608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd126609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd126610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=58;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=32337;
 end   
19'd126611: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=94;
   mapp<=46;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=33637;
 end   
19'd126612: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=54;
   mapp<=20;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=29854;
 end   
19'd126613: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=94;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd126614: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=13;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd126615: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=38;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd126616: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=98;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd126617: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd126618: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd126619: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd126761: begin  
rid<=1;
end
19'd126762: begin  
end
19'd126763: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd126764: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd126765: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd126766: begin  
rid<=0;
end
19'd126901: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=73;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3723;
 end   
19'd126902: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=19;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=4616;
 end   
19'd126903: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd127045: begin  
rid<=1;
end
19'd127046: begin  
end
19'd127047: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd127048: begin  
rid<=0;
end
19'd127201: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=99;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9083;
 end   
19'd127202: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=9;
   mapp<=46;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=14223;
 end   
19'd127203: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=56;
   mapp<=0;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8097;
 end   
19'd127204: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=43;
   mapp<=98;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=13976;
 end   
19'd127205: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=97;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=13132;
 end   
19'd127206: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd127207: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd127208: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd127209: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=64;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=26529;
 end   
19'd127210: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=54;
   mapp<=90;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=30235;
 end   
19'd127211: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=67;
   mapp<=74;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=23898;
 end   
19'd127212: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=30;
   mapp<=58;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=30040;
 end   
19'd127213: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=79;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=27831;
 end   
19'd127214: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd127215: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd127216: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd127217: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd127359: begin  
rid<=1;
end
19'd127360: begin  
end
19'd127361: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd127362: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd127363: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd127364: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd127365: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd127366: begin  
rid<=0;
end
19'd127501: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=76;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11667;
 end   
19'd127502: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=45;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11707;
 end   
19'd127503: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=53;
   mapp<=34;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9238;
 end   
19'd127504: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=35;
   mapp<=20;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=8354;
 end   
19'd127505: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=93;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=12328;
 end   
19'd127506: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=23;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7355;
 end   
19'd127507: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=40;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=7689;
 end   
19'd127508: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd127509: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd127510: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd127511: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=74;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=24377;
 end   
19'd127512: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=83;
   mapp<=26;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20893;
 end   
19'd127513: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=81;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=22050;
 end   
19'd127514: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=6;
   mapp<=12;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=18342;
 end   
19'd127515: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=80;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=25545;
 end   
19'd127516: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=26;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=19498;
 end   
19'd127517: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=59;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=23272;
 end   
19'd127518: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd127519: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd127520: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd127521: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd127663: begin  
rid<=1;
end
19'd127664: begin  
end
19'd127665: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd127666: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd127667: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd127668: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd127669: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd127670: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd127671: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd127672: begin  
rid<=0;
end
19'd127801: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=94;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10636;
 end   
19'd127802: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=30;
   mapp<=92;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9219;
 end   
19'd127803: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=30;
   mapp<=14;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6549;
 end   
19'd127804: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=14;
   mapp<=41;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=12740;
 end   
19'd127805: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=98;
   mapp<=5;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=13813;
 end   
19'd127806: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=39;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd127807: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=46;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd127808: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd127809: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=67;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd127810: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=92;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=20848;
 end   
19'd127811: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=14;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=17331;
 end   
19'd127812: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=87;
   mapp<=28;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=17405;
 end   
19'd127813: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=60;
   mapp<=30;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=20864;
 end   
19'd127814: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=14;
   mapp<=24;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=20267;
 end   
19'd127815: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=45;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd127816: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=64;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd127817: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=43;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd127818: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=19;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd127819: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd127961: begin  
rid<=1;
end
19'd127962: begin  
end
19'd127963: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd127964: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd127965: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd127966: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd127967: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd127968: begin  
rid<=0;
end
19'd128101: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=14;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=24570;
 end   
19'd128102: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=30;
   mapp<=63;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=26913;
 end   
19'd128103: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=79;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd128104: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=3;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd128105: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=99;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd128106: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=85;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd128107: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd128108: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=51;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd128109: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=54;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd128110: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=80;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd128111: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd128112: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=70;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=59404;
 end   
19'd128113: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=39;
   mapp<=8;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=59441;
 end   
19'd128114: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=52;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd128115: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=41;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd128116: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=44;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd128117: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=75;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd128118: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=72;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd128119: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=33;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd128120: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=94;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd128121: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=41;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd128122: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd128123: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd128265: begin  
rid<=1;
end
19'd128266: begin  
end
19'd128267: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd128268: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd128269: begin  
rid<=0;
end
19'd128401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=16;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=15011;
 end   
19'd128402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=97;
   mapp<=45;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=16042;
 end   
19'd128403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=88;
   mapp<=4;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=24292;
 end   
19'd128404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=16;
   mapp<=77;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=22631;
 end   
19'd128405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=56;
   mapp<=89;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=19910;
 end   
19'd128406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=28;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd128407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=29;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd128408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd128409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd128410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd128411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd128412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=46;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=41034;
 end   
19'd128413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=78;
   mapp<=46;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=37811;
 end   
19'd128414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=89;
   mapp<=87;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=46744;
 end   
19'd128415: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=98;
   mapp<=94;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=47368;
 end   
19'd128416: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=16;
   mapp<=14;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=37555;
 end   
19'd128417: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd128418: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=57;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd128419: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd128420: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd128421: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd128422: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd128423: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd128565: begin  
rid<=1;
end
19'd128566: begin  
end
19'd128567: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd128568: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd128569: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd128570: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd128571: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd128572: begin  
rid<=0;
end
19'd128701: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=25;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=15028;
 end   
19'd128702: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=84;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd128703: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=15;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd128704: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=52;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd128705: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=24;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd128706: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=18;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd128707: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=34;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=42575;
 end   
19'd128708: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=27;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd128709: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=25;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd128710: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=72;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd128711: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=88;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd128712: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=51;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd128713: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd128855: begin  
rid<=1;
end
19'd128856: begin  
end
19'd128857: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd128858: begin  
rid<=0;
end
19'd129001: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=70;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=18633;
 end   
19'd129002: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=11;
   mapp<=61;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12179;
 end   
19'd129003: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=33;
   mapp<=88;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=20159;
 end   
19'd129004: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=26;
   mapp<=39;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=18799;
 end   
19'd129005: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=52;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd129006: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=46;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd129007: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=21;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd129008: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=80;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd129009: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=36;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd129010: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=99;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=30117;
 end   
19'd129011: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=24;
   mapp<=45;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=25475;
 end   
19'd129012: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=29;
   mapp<=25;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=35581;
 end   
19'd129013: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=51;
   mapp<=23;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=31878;
 end   
19'd129014: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=28;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd129015: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=67;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd129016: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=98;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd129017: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=57;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd129018: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=41;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd129019: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd129161: begin  
rid<=1;
end
19'd129162: begin  
end
19'd129163: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd129164: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd129165: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd129166: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd129167: begin  
rid<=0;
end
19'd129301: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=15;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11394;
 end   
19'd129302: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=13;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8004;
 end   
19'd129303: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=49;
   mapp<=91;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8963;
 end   
19'd129304: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=24;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd129305: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=42;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd129306: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=54;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd129307: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=17;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd129308: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=40;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd129309: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=12;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd129310: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd129311: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd129312: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=18;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=36035;
 end   
19'd129313: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=20;
   mapp<=49;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=28411;
 end   
19'd129314: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=12;
   mapp<=28;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=33397;
 end   
19'd129315: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=97;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd129316: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=5;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd129317: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=46;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd129318: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=89;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd129319: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd129320: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=37;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd129321: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd129322: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd129323: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd129465: begin  
rid<=1;
end
19'd129466: begin  
end
19'd129467: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd129468: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd129469: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd129470: begin  
rid<=0;
end
19'd129601: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=28;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11118;
 end   
19'd129602: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=74;
   mapp<=92;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5923;
 end   
19'd129603: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=83;
   mapp<=17;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7173;
 end   
19'd129604: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=61;
   mapp<=3;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=10901;
 end   
19'd129605: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=30;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=11165;
 end   
19'd129606: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=65;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=13212;
 end   
19'd129607: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=52;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=14267;
 end   
19'd129608: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd129609: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd129610: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd129611: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=18;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17174;
 end   
19'd129612: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=5;
   mapp<=54;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=15679;
 end   
19'd129613: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=68;
   mapp<=24;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15095;
 end   
19'd129614: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=40;
   mapp<=98;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=20955;
 end   
19'd129615: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=50;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=18019;
 end   
19'd129616: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=90;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=19840;
 end   
19'd129617: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=48;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=17083;
 end   
19'd129618: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd129619: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd129620: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd129621: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd129763: begin  
rid<=1;
end
19'd129764: begin  
end
19'd129765: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd129766: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd129767: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd129768: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd129769: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd129770: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd129771: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd129772: begin  
rid<=0;
end
19'd129901: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=55;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1540;
 end   
19'd129902: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=35;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=990;
 end   
19'd129903: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=85;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2400;
 end   
19'd129904: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=29;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=1540;
 end   
19'd129905: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=54;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=990;
 end   
19'd129906: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=1;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=2400;
 end   
19'd129907: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd130049: begin  
rid<=1;
end
19'd130050: begin  
end
19'd130051: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd130052: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd130053: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd130054: begin  
rid<=0;
end
19'd130201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=10;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6768;
 end   
19'd130202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=47;
   mapp<=31;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7615;
 end   
19'd130203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=81;
   mapp<=61;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9236;
 end   
19'd130204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=55;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6677;
 end   
19'd130205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=74;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=9324;
 end   
19'd130206: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=38;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=4855;
 end   
19'd130207: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=88;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=4938;
 end   
19'd130208: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=11;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd130209: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=21;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd130210: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=97;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=9301;
 end   
19'd130211: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=31;
   mapp<=15;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8852;
 end   
19'd130212: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=43;
   mapp<=12;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=10932;
 end   
19'd130213: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=8;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=8743;
 end   
19'd130214: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=74;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=12167;
 end   
19'd130215: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=69;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=6931;
 end   
19'd130216: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=52;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=6778;
 end   
19'd130217: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd130218: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=64;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd130219: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd130361: begin  
rid<=1;
end
19'd130362: begin  
end
19'd130363: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd130364: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd130365: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd130366: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd130367: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd130368: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd130369: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd130370: begin  
rid<=0;
end
19'd130501: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=63;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10482;
 end   
19'd130502: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=76;
   mapp<=87;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8914;
 end   
19'd130503: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=1;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd130504: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=13;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd130505: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd130506: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=90;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=19179;
 end   
19'd130507: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=57;
   mapp<=88;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=13165;
 end   
19'd130508: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=18;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd130509: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=15;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd130510: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=17;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd130511: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd130653: begin  
rid<=1;
end
19'd130654: begin  
end
19'd130655: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd130656: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd130657: begin  
rid<=0;
end
19'd130801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=71;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6527;
 end   
19'd130802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=68;
   mapp<=49;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7039;
 end   
19'd130803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=81;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7144;
 end   
19'd130804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=71;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd130805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=86;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=9331;
 end   
19'd130806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=44;
   mapp<=52;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=9383;
 end   
19'd130807: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=40;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=8996;
 end   
19'd130808: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=31;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd130809: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd130951: begin  
rid<=1;
end
19'd130952: begin  
end
19'd130953: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd130954: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd130955: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd130956: begin  
rid<=0;
end
19'd131101: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=25;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=21199;
 end   
19'd131102: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=2;
   mapp<=59;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=19704;
 end   
19'd131103: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=20;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd131104: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=99;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd131105: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=34;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd131106: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=4;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd131107: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=69;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd131108: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=83;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd131109: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=68;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd131110: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=38;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd131111: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd131112: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=56;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=44032;
 end   
19'd131113: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=70;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=40171;
 end   
19'd131114: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=41;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd131115: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=39;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd131116: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=93;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd131117: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=96;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd131118: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=13;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd131119: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=31;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd131120: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=21;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd131121: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=72;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd131122: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd131123: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd131265: begin  
rid<=1;
end
19'd131266: begin  
end
19'd131267: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd131268: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd131269: begin  
rid<=0;
end
19'd131401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=25;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6460;
 end   
19'd131402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=75;
   mapp<=39;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10921;
 end   
19'd131403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=89;
   mapp<=15;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12715;
 end   
19'd131404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=99;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=14106;
 end   
19'd131405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=55;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=12877;
 end   
19'd131406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=84;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=13976;
 end   
19'd131407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd131408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd131409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=71;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=20680;
 end   
19'd131410: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=66;
   mapp<=94;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=24745;
 end   
19'd131411: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=35;
   mapp<=85;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=22354;
 end   
19'd131412: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=44;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=21175;
 end   
19'd131413: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=20;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=21382;
 end   
19'd131414: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=75;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=24167;
 end   
19'd131415: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd131416: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd131417: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd131559: begin  
rid<=1;
end
19'd131560: begin  
end
19'd131561: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd131562: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd131563: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd131564: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd131565: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd131566: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd131567: begin  
rid<=0;
end
19'd131701: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=39;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5453;
 end   
19'd131702: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=9;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5928;
 end   
19'd131703: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=57;
   mapp<=54;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7414;
 end   
19'd131704: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=2;
   mapp<=97;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7088;
 end   
19'd131705: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd131706: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd131707: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd131708: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=89;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=24183;
 end   
19'd131709: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=87;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18683;
 end   
19'd131710: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=97;
   mapp<=91;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=17101;
 end   
19'd131711: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=20;
   mapp<=2;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=18418;
 end   
19'd131712: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=67;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd131713: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=49;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd131714: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=26;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd131715: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd131857: begin  
rid<=1;
end
19'd131858: begin  
end
19'd131859: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd131860: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd131861: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd131862: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd131863: begin  
rid<=0;
end
19'd132001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=53;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=29286;
 end   
19'd132002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=48;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=24422;
 end   
19'd132003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=45;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd132004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=4;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd132005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=12;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd132006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=16;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd132007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=55;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd132008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=98;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd132009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=62;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd132010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=57;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd132011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd132012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=18;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=45679;
 end   
19'd132013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=18;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=38425;
 end   
19'd132014: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=29;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd132015: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=61;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd132016: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=32;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd132017: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=58;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd132018: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=46;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd132019: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=60;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd132020: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=43;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd132021: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=23;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd132022: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd132023: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd132165: begin  
rid<=1;
end
19'd132166: begin  
end
19'd132167: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd132168: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd132169: begin  
rid<=0;
end
19'd132301: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=75;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14487;
 end   
19'd132302: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=74;
   mapp<=31;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=13675;
 end   
19'd132303: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=16;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd132304: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=81;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd132305: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=57;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd132306: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=65;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd132307: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=43;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd132308: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=59;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd132309: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=50;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd132310: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=61;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=33604;
 end   
19'd132311: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=63;
   mapp<=78;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=29641;
 end   
19'd132312: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=55;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd132313: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=14;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd132314: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=50;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd132315: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=68;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd132316: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=26;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd132317: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=17;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd132318: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=85;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd132319: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd132461: begin  
rid<=1;
end
19'd132462: begin  
end
19'd132463: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd132464: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd132465: begin  
rid<=0;
end
19'd132601: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=2;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11058;
 end   
19'd132602: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=99;
   mapp<=12;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=20274;
 end   
19'd132603: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=17;
   mapp<=92;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=18122;
 end   
19'd132604: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=9;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd132605: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=52;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd132606: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=90;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd132607: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd132608: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=44;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd132609: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=87;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=29065;
 end   
19'd132610: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=77;
   mapp<=70;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=32921;
 end   
19'd132611: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=9;
   mapp<=3;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=29606;
 end   
19'd132612: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=63;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd132613: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=73;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd132614: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=31;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd132615: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=72;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd132616: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=86;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd132617: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd132759: begin  
rid<=1;
end
19'd132760: begin  
end
19'd132761: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd132762: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd132763: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd132764: begin  
rid<=0;
end
19'd132901: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=7;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=20515;
 end   
19'd132902: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=84;
   mapp<=63;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=29435;
 end   
19'd132903: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=44;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd132904: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=22;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd132905: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=73;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd132906: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=94;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd132907: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=73;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd132908: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=4;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd132909: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=59;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd132910: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=29;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd132911: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=62;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=45440;
 end   
19'd132912: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=92;
   mapp<=47;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=61276;
 end   
19'd132913: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=58;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd132914: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=98;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd132915: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=31;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd132916: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=79;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd132917: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=88;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd132918: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=73;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd132919: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=46;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd132920: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd132921: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd133063: begin  
rid<=1;
end
19'd133064: begin  
end
19'd133065: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd133066: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd133067: begin  
rid<=0;
end
19'd133201: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=41;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7840;
 end   
19'd133202: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=98;
   mapp<=80;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11816;
 end   
19'd133203: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=87;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7605;
 end   
19'd133204: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=41;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7689;
 end   
19'd133205: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd133206: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=8;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=11545;
 end   
19'd133207: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=41;
   mapp<=73;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12728;
 end   
19'd133208: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=8;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=8038;
 end   
19'd133209: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=9;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=9811;
 end   
19'd133210: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd133211: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd133353: begin  
rid<=1;
end
19'd133354: begin  
end
19'd133355: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd133356: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd133357: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd133358: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd133359: begin  
rid<=0;
end
19'd133501: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=35;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7602;
 end   
19'd133502: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=15;
   mapp<=4;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7584;
 end   
19'd133503: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=4;
   mapp<=36;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10491;
 end   
19'd133504: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=44;
   mapp<=67;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=8315;
 end   
19'd133505: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=50;
   mapp<=54;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5869;
 end   
19'd133506: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd133507: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd133508: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd133509: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd133510: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=73;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=25535;
 end   
19'd133511: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=89;
   mapp<=19;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=24103;
 end   
19'd133512: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=97;
   mapp<=81;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=27235;
 end   
19'd133513: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=38;
   mapp<=19;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=23700;
 end   
19'd133514: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=76;
   mapp<=48;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=24850;
 end   
19'd133515: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd133516: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd133517: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd133518: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd133519: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd133661: begin  
rid<=1;
end
19'd133662: begin  
end
19'd133663: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd133664: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd133665: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd133666: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd133667: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd133668: begin  
rid<=0;
end
19'd133801: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=89;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14541;
 end   
19'd133802: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=98;
   mapp<=29;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11993;
 end   
19'd133803: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=83;
   mapp<=50;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9290;
 end   
19'd133804: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=49;
   mapp<=36;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7106;
 end   
19'd133805: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=21;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5610;
 end   
19'd133806: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=39;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=8382;
 end   
19'd133807: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd133808: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd133809: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=84;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd133810: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=42;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=19093;
 end   
19'd133811: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=22;
   mapp<=22;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=16914;
 end   
19'd133812: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=16;
   mapp<=87;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=19536;
 end   
19'd133813: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=22;
   mapp<=93;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=23322;
 end   
19'd133814: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=25;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=22243;
 end   
19'd133815: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=79;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=24349;
 end   
19'd133816: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=91;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd133817: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=71;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd133818: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=71;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd133819: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd133961: begin  
rid<=1;
end
19'd133962: begin  
end
19'd133963: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd133964: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd133965: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd133966: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd133967: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd133968: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd133969: begin  
rid<=0;
end
19'd134101: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=67;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9080;
 end   
19'd134102: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=92;
   mapp<=62;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15392;
 end   
19'd134103: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=32;
   mapp<=83;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=16845;
 end   
19'd134104: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=8;
   mapp<=90;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=15520;
 end   
19'd134105: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=89;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=10623;
 end   
19'd134106: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=17;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=10297;
 end   
19'd134107: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=91;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=8477;
 end   
19'd134108: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=18;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=3812;
 end   
19'd134109: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd134110: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd134111: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd134112: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=36;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17757;
 end   
19'd134113: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=47;
   mapp<=98;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=30966;
 end   
19'd134114: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=23;
   mapp<=58;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=21780;
 end   
19'd134115: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=97;
   mapp<=13;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=28821;
 end   
19'd134116: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=93;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=17571;
 end   
19'd134117: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=1;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=16536;
 end   
19'd134118: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=87;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=14521;
 end   
19'd134119: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=16;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=12244;
 end   
19'd134120: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd134121: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd134122: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd134123: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd134265: begin  
rid<=1;
end
19'd134266: begin  
end
19'd134267: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd134268: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd134269: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd134270: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd134271: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd134272: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd134273: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd134274: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd134275: begin  
rid<=0;
end
19'd134401: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=48;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2512;
 end   
19'd134402: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=10;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3638;
 end   
19'd134403: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=44;
   mapp<=28;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2350;
 end   
19'd134404: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=15;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=2832;
 end   
19'd134405: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd134406: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd134407: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=44;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5740;
 end   
19'd134408: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=17;
   mapp<=4;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=7010;
 end   
19'd134409: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=68;
   mapp<=40;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=5555;
 end   
19'd134410: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=37;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6976;
 end   
19'd134411: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd134412: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd134413: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd134555: begin  
rid<=1;
end
19'd134556: begin  
end
19'd134557: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd134558: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd134559: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd134560: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd134561: begin  
rid<=0;
end
19'd134701: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=97;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8663;
 end   
19'd134702: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=46;
   mapp<=16;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4423;
 end   
19'd134703: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=53;
   mapp<=91;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9182;
 end   
19'd134704: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd134705: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=78;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd134706: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=28;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=18365;
 end   
19'd134707: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=24;
   mapp<=62;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18247;
 end   
19'd134708: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=81;
   mapp<=90;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=19623;
 end   
19'd134709: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd134710: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=25;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd134711: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd134853: begin  
rid<=1;
end
19'd134854: begin  
end
19'd134855: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd134856: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd134857: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd134858: begin  
rid<=0;
end
19'd135001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=67;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=15922;
 end   
19'd135002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=37;
   mapp<=96;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=17087;
 end   
19'd135003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=55;
   mapp<=62;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=19108;
 end   
19'd135004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=75;
   mapp<=63;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=18248;
 end   
19'd135005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=54;
   mapp<=35;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=18541;
 end   
19'd135006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=70;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=16797;
 end   
19'd135007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=63;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=16229;
 end   
19'd135008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=60;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd135009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=63;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd135010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd135011: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=94;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd135012: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=24;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=23980;
 end   
19'd135013: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=34;
   mapp<=18;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=25690;
 end   
19'd135014: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=6;
   mapp<=9;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=24014;
 end   
19'd135015: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=81;
   mapp<=64;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=25685;
 end   
19'd135016: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=90;
   mapp<=12;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=28446;
 end   
19'd135017: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=34;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=24571;
 end   
19'd135018: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=15;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=20298;
 end   
19'd135019: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd135020: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=80;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd135021: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=19;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd135022: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=26;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd135023: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd135165: begin  
rid<=1;
end
19'd135166: begin  
end
19'd135167: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd135168: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd135169: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd135170: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd135171: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd135172: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd135173: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd135174: begin  
rid<=0;
end
19'd135301: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=61;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3176;
 end   
19'd135302: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=22;
   mapp<=18;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1502;
 end   
19'd135303: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=6;
   mapp<=16;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=800;
 end   
19'd135304: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=26;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1852;
 end   
19'd135305: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=3;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1034;
 end   
19'd135306: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=39;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=2170;
 end   
19'd135307: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=10;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=1568;
 end   
19'd135308: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=14;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=2116;
 end   
19'd135309: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=51;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=4260;
 end   
19'd135310: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=32;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd135311: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=85;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd135312: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=2;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5647;
 end   
19'd135313: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=63;
   mapp<=1;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=7278;
 end   
19'd135314: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=64;
   mapp<=35;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=7588;
 end   
19'd135315: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=12;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=3285;
 end   
19'd135316: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=40;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=5700;
 end   
19'd135317: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=11;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=5861;
 end   
19'd135318: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=37;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=7589;
 end   
19'd135319: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=78;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=9939;
 end   
19'd135320: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=81;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=12883;
 end   
19'd135321: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd135322: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=51;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd135323: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd135465: begin  
rid<=1;
end
19'd135466: begin  
end
19'd135467: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd135468: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd135469: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd135470: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd135471: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd135472: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd135473: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd135474: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd135475: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd135476: begin  
rid<=0;
end
19'd135601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=88;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6851;
 end   
19'd135602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=75;
   mapp<=7;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6094;
 end   
19'd135603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=25;
   mapp<=49;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12109;
 end   
19'd135604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=7;
   mapp<=51;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=11071;
 end   
19'd135605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=28;
   mapp<=50;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=8350;
 end   
19'd135606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd135607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd135608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd135609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd135610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=6;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=27194;
 end   
19'd135611: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=16;
   mapp<=86;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=27259;
 end   
19'd135612: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=91;
   mapp<=73;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=30622;
 end   
19'd135613: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=51;
   mapp<=89;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=30710;
 end   
19'd135614: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=87;
   mapp<=85;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=27776;
 end   
19'd135615: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd135616: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd135617: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd135618: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd135619: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd135761: begin  
rid<=1;
end
19'd135762: begin  
end
19'd135763: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd135764: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd135765: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd135766: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd135767: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd135768: begin  
rid<=0;
end
19'd135901: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=25;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3855;
 end   
19'd135902: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=40;
   mapp<=52;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5110;
 end   
19'd135903: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=95;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3235;
 end   
19'd135904: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=21;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=595;
 end   
19'd135905: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=1;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3545;
 end   
19'd135906: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=87;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=3305;
 end   
19'd135907: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd135908: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=17;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7052;
 end   
19'd135909: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=55;
   mapp<=30;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8755;
 end   
19'd135910: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=57;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=7009;
 end   
19'd135911: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=51;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=1682;
 end   
19'd135912: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=4;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=7573;
 end   
19'd135913: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=72;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=5684;
 end   
19'd135914: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd135915: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd136057: begin  
rid<=1;
end
19'd136058: begin  
end
19'd136059: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd136060: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd136061: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd136062: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd136063: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd136064: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd136065: begin  
rid<=0;
end
19'd136201: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=78;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11866;
 end   
19'd136202: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=59;
   mapp<=98;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12728;
 end   
19'd136203: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=86;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11920;
 end   
19'd136204: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=88;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=8133;
 end   
19'd136205: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=21;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2327;
 end   
19'd136206: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=11;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=908;
 end   
19'd136207: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=1712;
 end   
19'd136208: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=28;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=2785;
 end   
19'd136209: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=9;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=2080;
 end   
19'd136210: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd136211: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=26;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16135;
 end   
19'd136212: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=49;
   mapp<=59;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=17594;
 end   
19'd136213: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=68;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15697;
 end   
19'd136214: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=41;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=10032;
 end   
19'd136215: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=17;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=5709;
 end   
19'd136216: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=60;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=5065;
 end   
19'd136217: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=53;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=5540;
 end   
19'd136218: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=50;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=8299;
 end   
19'd136219: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=86;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=4659;
 end   
19'd136220: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd136221: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd136363: begin  
rid<=1;
end
19'd136364: begin  
end
19'd136365: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd136366: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd136367: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd136368: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd136369: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd136370: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd136371: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd136372: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd136373: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd136374: begin  
rid<=0;
end
19'd136501: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=68;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12027;
 end   
19'd136502: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=8;
   mapp<=70;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12610;
 end   
19'd136503: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=59;
   mapp<=95;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=14513;
 end   
19'd136504: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=70;
   mapp<=22;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=10528;
 end   
19'd136505: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=53;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd136506: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=4;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd136507: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd136508: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd136509: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd136510: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=93;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=24292;
 end   
19'd136511: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=91;
   mapp<=54;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=22929;
 end   
19'd136512: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=40;
   mapp<=3;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=21124;
 end   
19'd136513: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=57;
   mapp<=1;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=19800;
 end   
19'd136514: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=17;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd136515: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=65;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd136516: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd136517: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd136518: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd136519: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd136661: begin  
rid<=1;
end
19'd136662: begin  
end
19'd136663: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd136664: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd136665: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd136666: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd136667: begin  
rid<=0;
end
19'd136801: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=23;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11205;
 end   
19'd136802: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=18;
   mapp<=88;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=16123;
 end   
19'd136803: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=87;
   mapp<=55;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12858;
 end   
19'd136804: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=96;
   mapp<=45;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5233;
 end   
19'd136805: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=7;
   mapp<=54;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=10820;
 end   
19'd136806: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=51;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=10936;
 end   
19'd136807: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=22;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=9679;
 end   
19'd136808: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=4;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd136809: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=90;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd136810: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=81;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd136811: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=10;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd136812: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=64;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=23993;
 end   
19'd136813: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=54;
   mapp<=17;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=27480;
 end   
19'd136814: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=93;
   mapp<=44;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=27621;
 end   
19'd136815: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=59;
   mapp<=12;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=16926;
 end   
19'd136816: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=57;
   mapp<=14;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=22308;
 end   
19'd136817: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=86;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=22599;
 end   
19'd136818: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=79;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=21768;
 end   
19'd136819: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=15;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd136820: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=56;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd136821: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=40;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd136822: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=82;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd136823: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd136965: begin  
rid<=1;
end
19'd136966: begin  
end
19'd136967: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd136968: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd136969: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd136970: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd136971: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd136972: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd136973: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd136974: begin  
rid<=0;
end
19'd137101: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=58;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=22800;
 end   
19'd137102: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=83;
   mapp<=82;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=13722;
 end   
19'd137103: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=52;
   mapp<=31;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=17482;
 end   
19'd137104: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=98;
   mapp<=90;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=11995;
 end   
19'd137105: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=7;
   mapp<=13;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=12425;
 end   
19'd137106: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=53;
   mapp<=31;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=14804;
 end   
19'd137107: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd137108: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd137109: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd137110: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd137111: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd137112: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=34;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=39514;
 end   
19'd137113: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=82;
   mapp<=22;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=31925;
 end   
19'd137114: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=31;
   mapp<=85;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=36706;
 end   
19'd137115: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=46;
   mapp<=84;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=29602;
 end   
19'd137116: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=70;
   mapp<=41;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=27461;
 end   
19'd137117: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=55;
   mapp<=55;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=25386;
 end   
19'd137118: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd137119: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd137120: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd137121: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd137122: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd137123: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd137265: begin  
rid<=1;
end
19'd137266: begin  
end
19'd137267: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd137268: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd137269: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd137270: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd137271: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd137272: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd137273: begin  
rid<=0;
end
19'd137401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=27;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7860;
 end   
19'd137402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=82;
   mapp<=60;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=13956;
 end   
19'd137403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=10;
   mapp<=78;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8380;
 end   
19'd137404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=87;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=12066;
 end   
19'd137405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=30;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd137406: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=42;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd137407: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=12;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=11861;
 end   
19'd137408: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=70;
   mapp<=53;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=16168;
 end   
19'd137409: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=15;
   mapp<=17;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=12681;
 end   
19'd137410: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=71;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=13918;
 end   
19'd137411: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=29;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd137412: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=6;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd137413: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd137555: begin  
rid<=1;
end
19'd137556: begin  
end
19'd137557: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd137558: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd137559: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd137560: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd137561: begin  
rid<=0;
end
19'd137701: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=4;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=20034;
 end   
19'd137702: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=45;
   mapp<=15;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=20213;
 end   
19'd137703: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=52;
   mapp<=67;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=20694;
 end   
19'd137704: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=81;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd137705: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=33;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd137706: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=50;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd137707: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=38;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd137708: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=72;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd137709: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=37;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd137710: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd137711: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd137712: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=29;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=39220;
 end   
19'd137713: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=95;
   mapp<=61;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=36784;
 end   
19'd137714: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=66;
   mapp<=56;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=31760;
 end   
19'd137715: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=25;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd137716: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=68;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd137717: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=25;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd137718: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=4;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd137719: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=44;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd137720: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=6;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd137721: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd137722: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd137723: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd137865: begin  
rid<=1;
end
19'd137866: begin  
end
19'd137867: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd137868: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd137869: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd137870: begin  
rid<=0;
end
19'd138001: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=97;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9506;
 end   
19'd138002: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=51;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4957;
 end   
19'd138003: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=34;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3318;
 end   
19'd138004: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=62;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6044;
 end   
19'd138005: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=34;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3338;
 end   
19'd138006: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=42;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=4124;
 end   
19'd138007: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=7;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=739;
 end   
19'd138008: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=89;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=8703;
 end   
19'd138009: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=27;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=10478;
 end   
19'd138010: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=89;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=7360;
 end   
19'd138011: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=44;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=4506;
 end   
19'd138012: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=51;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=7421;
 end   
19'd138013: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=64;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=5066;
 end   
19'd138014: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=73;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=6095;
 end   
19'd138015: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=79;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=2872;
 end   
19'd138016: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=55;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=10188;
 end   
19'd138017: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd138159: begin  
rid<=1;
end
19'd138160: begin  
end
19'd138161: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd138162: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd138163: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd138164: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd138165: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd138166: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd138167: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd138168: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd138169: begin  
rid<=0;
end
19'd138301: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=28;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4460;
 end   
19'd138302: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=15;
   mapp<=50;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6060;
 end   
19'd138303: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=35;
   mapp<=86;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4078;
 end   
19'd138304: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=96;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4943;
 end   
19'd138305: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=6;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2488;
 end   
19'd138306: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd138307: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd138308: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=65;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=10992;
 end   
19'd138309: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=3;
   mapp<=63;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=13133;
 end   
19'd138310: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=32;
   mapp<=54;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=8812;
 end   
19'd138311: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=88;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=12865;
 end   
19'd138312: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=30;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=4796;
 end   
19'd138313: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd138314: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd138315: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd138457: begin  
rid<=1;
end
19'd138458: begin  
end
19'd138459: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd138460: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd138461: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd138462: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd138463: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd138464: begin  
rid<=0;
end
19'd138601: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=20;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=15330;
 end   
19'd138602: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=88;
   mapp<=82;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8601;
 end   
19'd138603: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=12;
   mapp<=34;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10964;
 end   
19'd138604: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=41;
   mapp<=96;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=11241;
 end   
19'd138605: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=30;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd138606: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd138607: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd138608: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd138609: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=73;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=22089;
 end   
19'd138610: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=78;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18574;
 end   
19'd138611: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=74;
   mapp<=35;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=23973;
 end   
19'd138612: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=10;
   mapp<=78;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=25952;
 end   
19'd138613: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=19;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd138614: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd138615: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd138616: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd138617: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd138759: begin  
rid<=1;
end
19'd138760: begin  
end
19'd138761: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd138762: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd138763: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd138764: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd138765: begin  
rid<=0;
end
19'd138901: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=98;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1784;
 end   
19'd138902: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=48;
   mapp<=29;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1275;
 end   
19'd138903: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=37;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1821;
 end   
19'd138904: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=57;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1766;
 end   
19'd138905: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=52;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1553;
 end   
19'd138906: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=45;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=2985;
 end   
19'd138907: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=95;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=2557;
 end   
19'd138908: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=73;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=2537;
 end   
19'd138909: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=75;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd138910: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=82;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=6690;
 end   
19'd138911: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=33;
   mapp<=94;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=7641;
 end   
19'd138912: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=60;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=7841;
 end   
19'd138913: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=50;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=10856;
 end   
19'd138914: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=85;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=7559;
 end   
19'd138915: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=44;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=11755;
 end   
19'd138916: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=83;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=4947;
 end   
19'd138917: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=6;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=3703;
 end   
19'd138918: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=11;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd138919: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd139061: begin  
rid<=1;
end
19'd139062: begin  
end
19'd139063: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd139064: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd139065: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd139066: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd139067: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd139068: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd139069: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd139070: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd139071: begin  
rid<=0;
end
19'd139201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=94;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=15160;
 end   
19'd139202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=81;
   mapp<=92;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9306;
 end   
19'd139203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd139204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=18;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16911;
 end   
19'd139205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=13;
   mapp<=53;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=11300;
 end   
19'd139206: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd139207: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd139349: begin  
rid<=1;
end
19'd139350: begin  
end
19'd139351: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd139352: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd139353: begin  
rid<=0;
end
19'd139501: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=23;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=19580;
 end   
19'd139502: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=34;
   mapp<=64;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=19990;
 end   
19'd139503: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=39;
   mapp<=79;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=18847;
 end   
19'd139504: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=4;
   mapp<=94;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=18064;
 end   
19'd139505: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=75;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd139506: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=40;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd139507: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=34;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd139508: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=32;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd139509: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd139510: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=31;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd139511: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=98;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd139512: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=98;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=51945;
 end   
19'd139513: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=67;
   mapp<=69;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=50273;
 end   
19'd139514: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=81;
   mapp<=68;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=46155;
 end   
19'd139515: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=39;
   mapp<=82;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=49571;
 end   
19'd139516: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=91;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd139517: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=14;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd139518: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=82;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd139519: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=33;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd139520: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd139521: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=95;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd139522: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=99;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd139523: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd139665: begin  
rid<=1;
end
19'd139666: begin  
end
19'd139667: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd139668: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd139669: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd139670: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd139671: begin  
rid<=0;
end
19'd139801: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=62;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13081;
 end   
19'd139802: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=42;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=13027;
 end   
19'd139803: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=91;
   mapp<=72;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=14475;
 end   
19'd139804: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=83;
   mapp<=11;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=11914;
 end   
19'd139805: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=91;
   mapp<=16;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=9290;
 end   
19'd139806: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=45;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=10417;
 end   
19'd139807: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=28;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd139808: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=86;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd139809: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=53;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd139810: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=42;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd139811: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=81;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=30109;
 end   
19'd139812: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=60;
   mapp<=64;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=28802;
 end   
19'd139813: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=74;
   mapp<=33;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=30866;
 end   
19'd139814: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=51;
   mapp<=52;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=26273;
 end   
19'd139815: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=47;
   mapp<=24;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=23607;
 end   
19'd139816: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=73;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=24749;
 end   
19'd139817: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=59;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd139818: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd139819: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=18;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd139820: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=54;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd139821: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd139963: begin  
rid<=1;
end
19'd139964: begin  
end
19'd139965: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd139966: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd139967: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd139968: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd139969: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd139970: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd139971: begin  
rid<=0;
end
19'd140101: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7820;
 end   
19'd140102: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=1;
   mapp<=76;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7105;
 end   
19'd140103: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=63;
   mapp<=90;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7538;
 end   
19'd140104: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=34;
   mapp<=61;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3390;
 end   
19'd140105: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=93;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1844;
 end   
19'd140106: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=47;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=5494;
 end   
19'd140107: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=9;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=8630;
 end   
19'd140108: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=35;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=6658;
 end   
19'd140109: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd140110: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd140111: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd140112: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=85;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=18276;
 end   
19'd140113: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=85;
   mapp<=65;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20374;
 end   
19'd140114: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=8;
   mapp<=88;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=17710;
 end   
19'd140115: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=58;
   mapp<=4;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=8856;
 end   
19'd140116: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=4;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=9158;
 end   
19'd140117: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=40;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=16021;
 end   
19'd140118: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=77;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=21680;
 end   
19'd140119: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=51;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=12240;
 end   
19'd140120: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd140121: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd140122: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd140123: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd140265: begin  
rid<=1;
end
19'd140266: begin  
end
19'd140267: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd140268: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd140269: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd140270: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd140271: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd140272: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd140273: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd140274: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd140275: begin  
rid<=0;
end
19'd140401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=88;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12443;
 end   
19'd140402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=31;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=13362;
 end   
19'd140403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=10;
   mapp<=74;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=20737;
 end   
19'd140404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=70;
   mapp<=6;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=18623;
 end   
19'd140405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=49;
   mapp<=6;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=21767;
 end   
19'd140406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=65;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd140407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=72;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd140408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd140409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd140410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd140411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd140412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=38;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=26406;
 end   
19'd140413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=83;
   mapp<=99;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=25392;
 end   
19'd140414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=10;
   mapp<=30;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=34464;
 end   
19'd140415: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=27;
   mapp<=94;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=29803;
 end   
19'd140416: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=26;
   mapp<=16;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=33679;
 end   
19'd140417: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=24;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd140418: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=40;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd140419: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd140420: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd140421: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd140422: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd140423: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd140565: begin  
rid<=1;
end
19'd140566: begin  
end
19'd140567: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd140568: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd140569: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd140570: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd140571: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd140572: begin  
rid<=0;
end
19'd140701: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=79;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4941;
 end   
19'd140702: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=7;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2223;
 end   
19'd140703: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=45;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3675;
 end   
19'd140704: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=25;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4185;
 end   
19'd140705: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=67;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4433;
 end   
19'd140706: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=11;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=2299;
 end   
19'd140707: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=40;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=6300;
 end   
19'd140708: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=97;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd140709: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=26;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=10871;
 end   
19'd140710: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=68;
   mapp<=70;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=6473;
 end   
19'd140711: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=17;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=9340;
 end   
19'd140712: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=70;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=8385;
 end   
19'd140713: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=15;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=8118;
 end   
19'd140714: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=43;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=4234;
 end   
19'd140715: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=7840;
 end   
19'd140716: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=22;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd140717: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd140859: begin  
rid<=1;
end
19'd140860: begin  
end
19'd140861: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd140862: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd140863: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd140864: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd140865: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd140866: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd140867: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd140868: begin  
rid<=0;
end
19'd141001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=63;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6776;
 end   
19'd141002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=16;
   mapp<=28;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5979;
 end   
19'd141003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=35;
   mapp<=60;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7039;
 end   
19'd141004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=4;
   mapp<=67;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7655;
 end   
19'd141005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=18;
   mapp<=45;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5735;
 end   
19'd141006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=40;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6394;
 end   
19'd141007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=24;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=5120;
 end   
19'd141008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd141009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd141010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd141011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd141012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=13;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=20560;
 end   
19'd141013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=70;
   mapp<=8;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20294;
 end   
19'd141014: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=89;
   mapp<=94;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=18793;
 end   
19'd141015: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=49;
   mapp<=18;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=21200;
 end   
19'd141016: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=81;
   mapp<=47;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=19117;
 end   
19'd141017: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=46;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=21363;
 end   
19'd141018: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=35;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=21984;
 end   
19'd141019: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd141020: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd141021: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd141022: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd141023: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd141165: begin  
rid<=1;
end
19'd141166: begin  
end
19'd141167: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd141168: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd141169: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd141170: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd141171: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd141172: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd141173: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd141174: begin  
rid<=0;
end
19'd141301: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=6;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=108;
 end   
19'd141302: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=34;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=622;
 end   
19'd141303: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=81;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=1485;
 end   
19'd141304: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=22;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=996;
 end   
19'd141305: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd141447: begin  
rid<=1;
end
19'd141448: begin  
end
19'd141449: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd141450: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd141451: begin  
rid<=0;
end
19'd141601: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=24;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1752;
 end   
19'd141602: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=97;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7091;
 end   
19'd141603: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=87;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6371;
 end   
19'd141604: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=94;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6892;
 end   
19'd141605: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=48;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3544;
 end   
19'd141606: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=86;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6328;
 end   
19'd141607: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=14;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=1082;
 end   
19'd141608: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=94;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=6932;
 end   
19'd141609: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=41;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=2941;
 end   
19'd141610: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=81;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=9440;
 end   
19'd141611: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=23;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=7038;
 end   
19'd141612: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=62;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=8690;
 end   
19'd141613: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=44;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=4820;
 end   
19'd141614: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=59;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=8039;
 end   
19'd141615: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=29;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=1923;
 end   
19'd141616: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=48;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=8324;
 end   
19'd141617: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd141759: begin  
rid<=1;
end
19'd141760: begin  
end
19'd141761: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd141762: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd141763: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd141764: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd141765: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd141766: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd141767: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd141768: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd141769: begin  
rid<=0;
end
19'd141901: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=47;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2726;
 end   
19'd141902: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=21;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1228;
 end   
19'd141903: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=79;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4602;
 end   
19'd141904: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=1;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=88;
 end   
19'd141905: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=27;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1606;
 end   
19'd141906: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=27;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=1616;
 end   
19'd141907: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=52;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=3298;
 end   
19'd141908: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=93;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=2251;
 end   
19'd141909: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=39;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=5031;
 end   
19'd141910: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=35;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=473;
 end   
19'd141911: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=78;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=2464;
 end   
19'd141912: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=13;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=1759;
 end   
19'd141913: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd142055: begin  
rid<=1;
end
19'd142056: begin  
end
19'd142057: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd142058: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd142059: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd142060: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd142061: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd142062: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd142063: begin  
rid<=0;
end
19'd142201: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=51;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1636;
 end   
19'd142202: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=72;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1360;
 end   
19'd142203: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=52;
   mapp<=13;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6211;
 end   
19'd142204: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=6;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=11188;
 end   
19'd142205: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=98;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=11698;
 end   
19'd142206: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=73;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=5977;
 end   
19'd142207: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=27;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=3045;
 end   
19'd142208: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd142209: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd142210: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=81;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14203;
 end   
19'd142211: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=55;
   mapp<=66;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=15280;
 end   
19'd142212: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=96;
   mapp<=18;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=16142;
 end   
19'd142213: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=79;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=27248;
 end   
19'd142214: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=43;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=27329;
 end   
19'd142215: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=76;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=22458;
 end   
19'd142216: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=83;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=18060;
 end   
19'd142217: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd142218: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd142219: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd142361: begin  
rid<=1;
end
19'd142362: begin  
end
19'd142363: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd142364: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd142365: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd142366: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd142367: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd142368: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd142369: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd142370: begin  
rid<=0;
end
19'd142501: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=95;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12382;
 end   
19'd142502: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=26;
   mapp<=98;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=13706;
 end   
19'd142503: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=46;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd142504: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=98;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd142505: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=26;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd142506: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd142507: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=80;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=30496;
 end   
19'd142508: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=28;
   mapp<=63;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=28150;
 end   
19'd142509: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=7;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd142510: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=76;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd142511: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=59;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd142512: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=27;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd142513: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd142655: begin  
rid<=1;
end
19'd142656: begin  
end
19'd142657: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd142658: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd142659: begin  
rid<=0;
end
19'd142801: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=54;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4014;
 end   
19'd142802: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=41;
   mapp<=90;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7207;
 end   
19'd142803: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=57;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5107;
 end   
19'd142804: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=49;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5710;
 end   
19'd142805: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd142806: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=85;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12127;
 end   
19'd142807: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=59;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=17351;
 end   
19'd142808: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=61;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=11295;
 end   
19'd142809: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=17;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=12760;
 end   
19'd142810: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd142811: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd142953: begin  
rid<=1;
end
19'd142954: begin  
end
19'd142955: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd142956: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd142957: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd142958: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd142959: begin  
rid<=0;
end
19'd143101: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=75;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=20349;
 end   
19'd143102: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=16;
   mapp<=16;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=22302;
 end   
19'd143103: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=45;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd143104: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=71;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd143105: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=62;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd143106: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=45;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd143107: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=30;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd143108: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=80;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd143109: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd143110: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=78;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=53324;
 end   
19'd143111: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=19;
   mapp<=98;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=57814;
 end   
19'd143112: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=96;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd143113: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=28;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd143114: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=89;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd143115: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=77;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd143116: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=56;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd143117: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=83;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd143118: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd143119: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd143261: begin  
rid<=1;
end
19'd143262: begin  
end
19'd143263: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd143264: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd143265: begin  
rid<=0;
end
19'd143401: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=45;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=18445;
 end   
19'd143402: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=48;
   mapp<=79;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=21713;
 end   
19'd143403: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=65;
   mapp<=98;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=19172;
 end   
19'd143404: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=67;
   mapp<=57;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=16729;
 end   
19'd143405: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=21;
   mapp<=69;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=18509;
 end   
19'd143406: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=81;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=16617;
 end   
19'd143407: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=41;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=19926;
 end   
19'd143408: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=4;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd143409: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=93;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd143410: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=32;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd143411: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=85;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd143412: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=91;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=38721;
 end   
19'd143413: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=67;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=41586;
 end   
19'd143414: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=6;
   mapp<=88;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=38226;
 end   
19'd143415: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=68;
   mapp<=81;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=40719;
 end   
19'd143416: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=92;
   mapp<=1;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=44493;
 end   
19'd143417: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=50;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=43141;
 end   
19'd143418: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=62;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=44688;
 end   
19'd143419: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=96;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd143420: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=98;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd143421: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=22;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd143422: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd143423: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd143565: begin  
rid<=1;
end
19'd143566: begin  
end
19'd143567: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd143568: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd143569: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd143570: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd143571: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd143572: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd143573: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd143574: begin  
rid<=0;
end
19'd143701: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=90;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4314;
 end   
19'd143702: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=39;
   mapp<=64;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5725;
 end   
19'd143703: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=18;
   mapp<=66;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5692;
 end   
19'd143704: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=65;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6383;
 end   
19'd143705: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=21;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=10477;
 end   
19'd143706: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=69;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=10057;
 end   
19'd143707: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=89;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=9609;
 end   
19'd143708: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=58;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=10944;
 end   
19'd143709: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=79;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=7795;
 end   
19'd143710: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=82;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd143711: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=29;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd143712: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=76;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=13852;
 end   
19'd143713: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=97;
   mapp<=90;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12503;
 end   
19'd143714: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=63;
   mapp<=8;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=14052;
 end   
19'd143715: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=90;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=7065;
 end   
19'd143716: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=1;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=13323;
 end   
19'd143717: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=29;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=13159;
 end   
19'd143718: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=29;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=14651;
 end   
19'd143719: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=47;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=19210;
 end   
19'd143720: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=87;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=10957;
 end   
19'd143721: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=31;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd143722: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=3;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd143723: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd143865: begin  
rid<=1;
end
19'd143866: begin  
end
19'd143867: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd143868: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd143869: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd143870: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd143871: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd143872: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd143873: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd143874: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd143875: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd143876: begin  
rid<=0;
end
19'd144001: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=69;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8095;
 end   
19'd144002: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=22;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd144003: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=64;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17621;
 end   
19'd144004: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=74;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd144005: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd144147: begin  
rid<=1;
end
19'd144148: begin  
end
19'd144149: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd144150: begin  
rid<=0;
end
19'd144301: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=39;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16220;
 end   
19'd144302: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=88;
   mapp<=86;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=17288;
 end   
19'd144303: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=65;
   mapp<=67;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=17693;
 end   
19'd144304: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=78;
   mapp<=5;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=15996;
 end   
19'd144305: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=98;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd144306: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=18;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd144307: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=6;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd144308: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd144309: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=24;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=21775;
 end   
19'd144310: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=33;
   mapp<=36;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=25039;
 end   
19'd144311: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=59;
   mapp<=61;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=22002;
 end   
19'd144312: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=56;
   mapp<=0;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=25385;
 end   
19'd144313: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=32;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd144314: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=99;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd144315: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=5;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd144316: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=94;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd144317: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd144459: begin  
rid<=1;
end
19'd144460: begin  
end
19'd144461: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd144462: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd144463: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd144464: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd144465: begin  
rid<=0;
end
19'd144601: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=54;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1782;
 end   
19'd144602: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5248;
 end   
19'd144603: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=92;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4988;
 end   
19'd144604: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=56;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3054;
 end   
19'd144605: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=85;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4630;
 end   
19'd144606: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=51;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=2804;
 end   
19'd144607: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=30;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=1680;
 end   
19'd144608: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=24;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=1366;
 end   
19'd144609: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=38;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=4784;
 end   
19'd144610: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=7984;
 end   
19'd144611: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=18;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=5672;
 end   
19'd144612: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=94;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6626;
 end   
19'd144613: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=47;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=6416;
 end   
19'd144614: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=23;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=3678;
 end   
19'd144615: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=36;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=3048;
 end   
19'd144616: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=72;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=4102;
 end   
19'd144617: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd144759: begin  
rid<=1;
end
19'd144760: begin  
end
19'd144761: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd144762: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd144763: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd144764: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd144765: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd144766: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd144767: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd144768: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd144769: begin  
rid<=0;
end
19'd144901: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=76;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9964;
 end   
19'd144902: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=56;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9602;
 end   
19'd144903: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=79;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7368;
 end   
19'd144904: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=24;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5494;
 end   
19'd144905: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=65;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6492;
 end   
19'd144906: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=27;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=4174;
 end   
19'd144907: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=37;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=4552;
 end   
19'd144908: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=30;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=7446;
 end   
19'd144909: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=91;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=9740;
 end   
19'd144910: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=49;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=5774;
 end   
19'd144911: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd144912: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=8;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=15864;
 end   
19'd144913: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=62;
   mapp<=90;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12554;
 end   
19'd144914: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=36;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=11376;
 end   
19'd144915: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=60;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=10748;
 end   
19'd144916: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=77;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=8782;
 end   
19'd144917: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=27;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=7924;
 end   
19'd144918: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=57;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=5442;
 end   
19'd144919: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=7;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=9734;
 end   
19'd144920: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=36;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=13004;
 end   
19'd144921: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=48;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=9940;
 end   
19'd144922: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd144923: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd145065: begin  
rid<=1;
end
19'd145066: begin  
end
19'd145067: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd145068: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd145069: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd145070: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd145071: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd145072: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd145073: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd145074: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd145075: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd145076: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd145077: begin  
rid<=0;
end
19'd145201: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=19;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9858;
 end   
19'd145202: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=19;
   mapp<=88;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12581;
 end   
19'd145203: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=98;
   mapp<=13;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11531;
 end   
19'd145204: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=66;
   mapp<=18;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=9667;
 end   
19'd145205: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=50;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd145206: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=18;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd145207: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=14;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd145208: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=56;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd145209: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd145210: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd145211: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd145212: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=77;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=33071;
 end   
19'd145213: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=81;
   mapp<=44;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=43776;
 end   
19'd145214: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=94;
   mapp<=63;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=39454;
 end   
19'd145215: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=57;
   mapp<=51;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=38700;
 end   
19'd145216: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=72;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd145217: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=71;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd145218: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=17;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd145219: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=94;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd145220: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd145221: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd145222: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd145223: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd145365: begin  
rid<=1;
end
19'd145366: begin  
end
19'd145367: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd145368: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd145369: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd145370: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd145371: begin  
rid<=0;
end
19'd145501: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=3;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7446;
 end   
19'd145502: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=88;
   mapp<=63;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6797;
 end   
19'd145503: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=49;
   mapp<=36;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8052;
 end   
19'd145504: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=70;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4682;
 end   
19'd145505: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=36;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4984;
 end   
19'd145506: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=26;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=8379;
 end   
19'd145507: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd145508: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd145509: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=85;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16144;
 end   
19'd145510: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=61;
   mapp<=43;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=14538;
 end   
19'd145511: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=28;
   mapp<=50;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=17275;
 end   
19'd145512: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=37;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=14640;
 end   
19'd145513: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=97;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=16385;
 end   
19'd145514: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=32;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=16074;
 end   
19'd145515: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd145516: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd145517: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd145659: begin  
rid<=1;
end
19'd145660: begin  
end
19'd145661: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd145662: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd145663: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd145664: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd145665: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd145666: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd145667: begin  
rid<=0;
end
19'd145801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=80;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=360;
 end   
19'd145802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=4;
   mapp<=10;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=566;
 end   
19'd145803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=54;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=456;
 end   
19'd145804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=22;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=898;
 end   
19'd145805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=78;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=822;
 end   
19'd145806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=47;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=268;
 end   
19'd145807: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=3;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=1062;
 end   
19'd145808: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=99;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=736;
 end   
19'd145809: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=27;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=538;
 end   
19'd145810: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=35;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd145811: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=75;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=11826;
 end   
19'd145812: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=62;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8440;
 end   
19'd145813: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=34;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=11038;
 end   
19'd145814: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=86;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=8736;
 end   
19'd145815: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=14;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=11093;
 end   
19'd145816: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=99;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=9094;
 end   
19'd145817: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=14;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=4079;
 end   
19'd145818: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=21;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=8377;
 end   
19'd145819: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=65;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=5943;
 end   
19'd145820: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=5;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd145821: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd145963: begin  
rid<=1;
end
19'd145964: begin  
end
19'd145965: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd145966: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd145967: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd145968: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd145969: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd145970: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd145971: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd145972: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd145973: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd145974: begin  
rid<=0;
end
19'd146101: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=2;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3416;
 end   
19'd146102: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=8;
   mapp<=38;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4107;
 end   
19'd146103: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd146104: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=33;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd146105: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=0;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd146106: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=8;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=19710;
 end   
19'd146107: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=80;
   mapp<=42;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18895;
 end   
19'd146108: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=80;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd146109: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=82;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd146110: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=0;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd146111: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd146253: begin  
rid<=1;
end
19'd146254: begin  
end
19'd146255: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd146256: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd146257: begin  
rid<=0;
end
19'd146401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=28;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4169;
 end   
19'd146402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=57;
   mapp<=25;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2819;
 end   
19'd146403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=37;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6243;
 end   
19'd146404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=91;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6283;
 end   
19'd146405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=65;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4311;
 end   
19'd146406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=43;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=3363;
 end   
19'd146407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=37;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=6625;
 end   
19'd146408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd146409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=34;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=6305;
 end   
19'd146410: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=6;
   mapp<=16;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=3777;
 end   
19'd146411: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=69;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=8955;
 end   
19'd146412: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=61;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=8771;
 end   
19'd146413: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=69;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=7041;
 end   
19'd146414: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=64;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=5539;
 end   
19'd146415: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=7027;
 end   
19'd146416: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd146417: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd146559: begin  
rid<=1;
end
19'd146560: begin  
end
19'd146561: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd146562: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd146563: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd146564: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd146565: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd146566: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd146567: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd146568: begin  
rid<=0;
end
19'd146701: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=33;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2805;
 end   
19'd146702: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=16;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=538;
 end   
19'd146703: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=50;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1670;
 end   
19'd146704: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=67;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=2241;
 end   
19'd146705: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=25;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=865;
 end   
19'd146706: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=4;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=182;
 end   
19'd146707: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=76;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=10025;
 end   
19'd146708: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=20;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=2058;
 end   
19'd146709: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=77;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=7522;
 end   
19'd146710: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=90;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=9081;
 end   
19'd146711: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=71;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=6261;
 end   
19'd146712: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=6;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=638;
 end   
19'd146713: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd146855: begin  
rid<=1;
end
19'd146856: begin  
end
19'd146857: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd146858: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd146859: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd146860: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd146861: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd146862: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd146863: begin  
rid<=0;
end
19'd147001: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=61;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=732;
 end   
19'd147002: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=74;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4524;
 end   
19'd147003: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=97;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5937;
 end   
19'd147004: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=3;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=213;
 end   
19'd147005: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=80;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5612;
 end   
19'd147006: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=10684;
 end   
19'd147007: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=10;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=6737;
 end   
19'd147008: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=84;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6933;
 end   
19'd147009: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd147151: begin  
rid<=1;
end
19'd147152: begin  
end
19'd147153: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd147154: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd147155: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd147156: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd147157: begin  
rid<=0;
end
19'd147301: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=7;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=560;
 end   
19'd147302: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=0;
   mapp<=30;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=220;
 end   
19'd147303: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=74;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=1966;
 end   
19'd147304: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=0;
   mapp<=13;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=1182;
 end   
19'd147305: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd147447: begin  
rid<=1;
end
19'd147448: begin  
end
19'd147449: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd147450: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd147451: begin  
rid<=0;
end
19'd147601: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=42;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7000;
 end   
19'd147602: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=56;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3146;
 end   
19'd147603: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd147604: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=6;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7648;
 end   
19'd147605: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=72;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8558;
 end   
19'd147606: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd147607: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd147749: begin  
rid<=1;
end
19'd147750: begin  
end
19'd147751: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd147752: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd147753: begin  
rid<=0;
end
19'd147901: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=15;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12547;
 end   
19'd147902: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=45;
   mapp<=55;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=14040;
 end   
19'd147903: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=97;
   mapp<=52;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12600;
 end   
19'd147904: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=61;
   mapp<=54;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=15598;
 end   
19'd147905: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=84;
   mapp<=11;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=18817;
 end   
19'd147906: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=59;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=19185;
 end   
19'd147907: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd147908: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd147909: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd147910: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd147911: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd147912: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=5;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=20437;
 end   
19'd147913: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=62;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=22690;
 end   
19'd147914: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=50;
   mapp<=82;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=21100;
 end   
19'd147915: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=59;
   mapp<=43;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=23837;
 end   
19'd147916: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=4;
   mapp<=82;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=26864;
 end   
19'd147917: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=16;
   mapp<=50;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=26285;
 end   
19'd147918: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd147919: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd147920: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd147921: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd147922: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd147923: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd148065: begin  
rid<=1;
end
19'd148066: begin  
end
19'd148067: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd148068: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd148069: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd148070: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd148071: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd148072: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd148073: begin  
rid<=0;
end
19'd148201: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=59;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=118;
 end   
19'd148202: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=31;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1839;
 end   
19'd148203: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=31;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1849;
 end   
19'd148204: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=3;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=207;
 end   
19'd148205: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=15;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=925;
 end   
19'd148206: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=97;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7975;
 end   
19'd148207: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=81;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=9696;
 end   
19'd148208: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=32;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=4953;
 end   
19'd148209: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=24;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=2535;
 end   
19'd148210: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=95;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=10140;
 end   
19'd148211: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd148353: begin  
rid<=1;
end
19'd148354: begin  
end
19'd148355: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd148356: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd148357: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd148358: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd148359: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd148360: begin  
rid<=0;
end
19'd148501: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=82;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5904;
 end   
19'd148502: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=56;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4042;
 end   
19'd148503: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=82;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5924;
 end   
19'd148504: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=93;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6726;
 end   
19'd148505: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=55;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8489;
 end   
19'd148506: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=28;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=5358;
 end   
19'd148507: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=43;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=7945;
 end   
19'd148508: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=62;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=9640;
 end   
19'd148509: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd148651: begin  
rid<=1;
end
19'd148652: begin  
end
19'd148653: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd148654: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd148655: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd148656: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd148657: begin  
rid<=0;
end
19'd148801: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=74;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14694;
 end   
19'd148802: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=64;
   mapp<=71;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=14553;
 end   
19'd148803: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=47;
   mapp<=86;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12015;
 end   
19'd148804: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=8;
   mapp<=79;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=8065;
 end   
19'd148805: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=9;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6896;
 end   
19'd148806: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=19;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=11715;
 end   
19'd148807: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd148808: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd148809: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd148810: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=5;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=25583;
 end   
19'd148811: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=84;
   mapp<=46;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=24796;
 end   
19'd148812: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=59;
   mapp<=50;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=21175;
 end   
19'd148813: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=80;
   mapp<=47;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=15978;
 end   
19'd148814: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=38;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=14011;
 end   
19'd148815: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=34;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=20461;
 end   
19'd148816: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd148817: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd148818: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd148819: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd148961: begin  
rid<=1;
end
19'd148962: begin  
end
19'd148963: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd148964: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd148965: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd148966: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd148967: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd148968: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd148969: begin  
rid<=0;
end
19'd149101: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=44;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=17493;
 end   
19'd149102: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=65;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=23173;
 end   
19'd149103: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=87;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=23946;
 end   
19'd149104: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=53;
   mapp<=87;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=22831;
 end   
19'd149105: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=74;
   mapp<=55;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=24351;
 end   
19'd149106: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=48;
   mapp<=83;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=22600;
 end   
19'd149107: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=93;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd149108: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=63;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd149109: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=18;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd149110: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=61;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd149111: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=68;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd149112: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=39;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=23206;
 end   
19'd149113: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=18;
   mapp<=63;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=32042;
 end   
19'd149114: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=28;
   mapp<=8;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=30505;
 end   
19'd149115: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=7;
   mapp<=48;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=29245;
 end   
19'd149116: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=67;
   mapp<=35;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=35330;
 end   
19'd149117: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=93;
   mapp<=5;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=28963;
 end   
19'd149118: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=4;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd149119: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=22;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd149120: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=54;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd149121: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=13;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd149122: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=1;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd149123: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd149265: begin  
rid<=1;
end
19'd149266: begin  
end
19'd149267: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd149268: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd149269: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd149270: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd149271: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd149272: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd149273: begin  
rid<=0;
end
19'd149401: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=84;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=840;
 end   
19'd149402: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=79;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6646;
 end   
19'd149403: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=42;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3548;
 end   
19'd149404: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=9;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=786;
 end   
19'd149405: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=75;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=3240;
 end   
19'd149406: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12871;
 end   
19'd149407: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=57;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=7823;
 end   
19'd149408: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=2;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=936;
 end   
19'd149409: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd149551: begin  
rid<=1;
end
19'd149552: begin  
end
19'd149553: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd149554: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd149555: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd149556: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd149557: begin  
rid<=0;
end
19'd149701: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=63;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3478;
 end   
19'd149702: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=17;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd149703: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=80;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5558;
 end   
19'd149704: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=72;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd149705: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd149847: begin  
rid<=1;
end
19'd149848: begin  
end
19'd149849: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd149850: begin  
rid<=0;
end
19'd150001: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=75;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3942;
 end   
19'd150002: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=81;
   mapp<=7;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5557;
 end   
19'd150003: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=62;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6776;
 end   
19'd150004: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd150005: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=10;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8738;
 end   
19'd150006: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=64;
   mapp<=69;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12135;
 end   
19'd150007: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=92;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=13328;
 end   
19'd150008: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd150009: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd150151: begin  
rid<=1;
end
19'd150152: begin  
end
19'd150153: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd150154: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd150155: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd150156: begin  
rid<=0;
end
19'd150301: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=71;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7266;
 end   
19'd150302: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=9;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=649;
 end   
19'd150303: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=25;
   mapp<=89;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7580;
 end   
19'd150304: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6883;
 end   
19'd150305: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=65;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=11597;
 end   
19'd150306: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=77;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd150307: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=78;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd150308: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=94;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=13102;
 end   
19'd150309: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=2;
   mapp<=26;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=1449;
 end   
19'd150310: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=25;
   mapp<=2;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=9553;
 end   
19'd150311: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=14;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=8975;
 end   
19'd150312: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=42;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=16059;
 end   
19'd150313: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=73;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd150314: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=1;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd150315: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd150457: begin  
rid<=1;
end
19'd150458: begin  
end
19'd150459: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd150460: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd150461: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd150462: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd150463: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd150464: begin  
rid<=0;
end
19'd150601: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=49;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5178;
 end   
19'd150602: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=29;
   mapp<=3;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2564;
 end   
19'd150603: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=59;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd150604: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd150605: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=61;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=15445;
 end   
19'd150606: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=96;
   mapp<=49;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12021;
 end   
19'd150607: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=3;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd150608: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd150609: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd150751: begin  
rid<=1;
end
19'd150752: begin  
end
19'd150753: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd150754: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd150755: begin  
rid<=0;
end
19'd150901: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=3;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=141;
 end   
19'd150902: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=94;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4428;
 end   
19'd150903: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=27;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1289;
 end   
19'd150904: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=74;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3508;
 end   
19'd150905: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=34;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1638;
 end   
19'd150906: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=91;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=4327;
 end   
19'd150907: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=59;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=2833;
 end   
19'd150908: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=5;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=305;
 end   
19'd150909: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=31;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=1537;
 end   
19'd150910: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=63;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5622;
 end   
19'd150911: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=13;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=5559;
 end   
19'd150912: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=5;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=1724;
 end   
19'd150913: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=74;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=9946;
 end   
19'd150914: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=23;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=3639;
 end   
19'd150915: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=85;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=11722;
 end   
19'd150916: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=51;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=7270;
 end   
19'd150917: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=98;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=8831;
 end   
19'd150918: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=47;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=5626;
 end   
19'd150919: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd151061: begin  
rid<=1;
end
19'd151062: begin  
end
19'd151063: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd151064: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd151065: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd151066: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd151067: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd151068: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd151069: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd151070: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd151071: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd151072: begin  
rid<=0;
end
19'd151201: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=50;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5490;
 end   
19'd151202: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=14;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd151203: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=80;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=13458;
 end   
19'd151204: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=16;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd151205: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd151347: begin  
rid<=1;
end
19'd151348: begin  
end
19'd151349: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd151350: begin  
rid<=0;
end
19'd151501: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=77;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=17767;
 end   
19'd151502: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=26;
   mapp<=31;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=17927;
 end   
19'd151503: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=62;
   mapp<=88;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=22649;
 end   
19'd151504: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=64;
   mapp<=8;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=13023;
 end   
19'd151505: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=67;
   mapp<=59;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=22226;
 end   
19'd151506: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=88;
   mapp<=38;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=23475;
 end   
19'd151507: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd151508: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd151509: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd151510: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd151511: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd151512: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=16;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=24879;
 end   
19'd151513: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=3;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=24203;
 end   
19'd151514: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=12;
   mapp<=92;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=27555;
 end   
19'd151515: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=74;
   mapp<=36;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=17298;
 end   
19'd151516: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=32;
   mapp<=51;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=30220;
 end   
19'd151517: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=26;
   mapp<=18;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=32124;
 end   
19'd151518: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd151519: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd151520: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd151521: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd151522: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd151523: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd151665: begin  
rid<=1;
end
19'd151666: begin  
end
19'd151667: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd151668: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd151669: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd151670: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd151671: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd151672: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd151673: begin  
rid<=0;
end
19'd151801: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=22;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1628;
 end   
19'd151802: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=53;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3932;
 end   
19'd151803: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=50;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3720;
 end   
19'd151804: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=30;
 end   
19'd151805: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=8;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=632;
 end   
19'd151806: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=24;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=1826;
 end   
19'd151807: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=3;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=282;
 end   
19'd151808: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=8;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=662;
 end   
19'd151809: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=77;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=5778;
 end   
19'd151810: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=27;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=2088;
 end   
19'd151811: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=21;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=3224;
 end   
19'd151812: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=91;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=10848;
 end   
19'd151813: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=91;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=10636;
 end   
19'd151814: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=65;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=4970;
 end   
19'd151815: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=49;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=4356;
 end   
19'd151816: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=36;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=4562;
 end   
19'd151817: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=7;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=814;
 end   
19'd151818: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=46;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=4158;
 end   
19'd151819: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=36;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=8514;
 end   
19'd151820: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=26;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=4064;
 end   
19'd151821: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd151963: begin  
rid<=1;
end
19'd151964: begin  
end
19'd151965: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd151966: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd151967: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd151968: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd151969: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd151970: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd151971: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd151972: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd151973: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd151974: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd151975: begin  
rid<=0;
end
19'd152101: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=11;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=15438;
 end   
19'd152102: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=25;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd152103: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=98;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd152104: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=40;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd152105: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=86;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd152106: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=83;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd152107: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=25;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd152108: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=99;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd152109: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=13;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=35554;
 end   
19'd152110: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=52;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd152111: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=34;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd152112: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=54;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd152113: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=32;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd152114: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=1;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd152115: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=31;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd152116: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=77;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd152117: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd152259: begin  
rid<=1;
end
19'd152260: begin  
end
19'd152261: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd152262: begin  
rid<=0;
end
19'd152401: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=80;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10044;
 end   
19'd152402: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=4;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=13079;
 end   
19'd152403: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=62;
   mapp<=79;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=13681;
 end   
19'd152404: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=4;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd152405: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=55;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd152406: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=35;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd152407: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=80;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd152408: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=82;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd152409: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=71;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd152410: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=95;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=29156;
 end   
19'd152411: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=10;
   mapp<=70;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=29272;
 end   
19'd152412: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=95;
   mapp<=64;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=29270;
 end   
19'd152413: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=5;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd152414: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=64;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd152415: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=56;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd152416: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=71;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd152417: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=11;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd152418: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=1;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd152419: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd152561: begin  
rid<=1;
end
19'd152562: begin  
end
19'd152563: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd152564: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd152565: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd152566: begin  
rid<=0;
end
19'd152701: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9727;
 end   
19'd152702: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=30;
   mapp<=51;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11091;
 end   
19'd152703: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=15;
   mapp<=60;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=13510;
 end   
19'd152704: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=10;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd152705: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=61;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd152706: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=78;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd152707: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=47;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd152708: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=42;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd152709: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd152710: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd152711: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=7;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=27612;
 end   
19'd152712: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=35;
   mapp<=20;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=27666;
 end   
19'd152713: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=20;
   mapp<=62;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=28204;
 end   
19'd152714: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=37;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd152715: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=42;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd152716: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=52;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd152717: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=82;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd152718: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=78;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd152719: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd152720: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd152721: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd152863: begin  
rid<=1;
end
19'd152864: begin  
end
19'd152865: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd152866: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd152867: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd152868: begin  
rid<=0;
end
19'd153001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=1;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7592;
 end   
19'd153002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd153003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=23;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd153004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=5;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd153005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=72;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd153006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=61;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=26611;
 end   
19'd153007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=86;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd153008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=69;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd153009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=93;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd153010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=24;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd153011: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd153153: begin  
rid<=1;
end
19'd153154: begin  
end
19'd153155: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd153156: begin  
rid<=0;
end
19'd153301: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=46;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7090;
 end   
19'd153302: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=32;
   mapp<=85;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8745;
 end   
19'd153303: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=67;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12845;
 end   
19'd153304: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=76;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7420;
 end   
19'd153305: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=2;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6775;
 end   
19'd153306: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=77;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=15780;
 end   
19'd153307: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=99;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=15755;
 end   
19'd153308: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=74;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=9735;
 end   
19'd153309: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=31;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=11440;
 end   
19'd153310: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=99;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=9750;
 end   
19'd153311: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=3;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd153312: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=42;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=13032;
 end   
19'd153313: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=50;
   mapp<=76;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18743;
 end   
19'd153314: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=98;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=19971;
 end   
19'd153315: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=28;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=14016;
 end   
19'd153316: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=68;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=13967;
 end   
19'd153317: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=49;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=22535;
 end   
19'd153318: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=56;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=24159;
 end   
19'd153319: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=73;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=18626;
 end   
19'd153320: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=68;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=18404;
 end   
19'd153321: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=46;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=13844;
 end   
19'd153322: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd153323: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd153465: begin  
rid<=1;
end
19'd153466: begin  
end
19'd153467: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd153468: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd153469: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd153470: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd153471: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd153472: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd153473: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd153474: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd153475: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd153476: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd153477: begin  
rid<=0;
end
19'd153601: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=17;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=765;
 end   
19'd153602: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1591;
 end   
19'd153603: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=44;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=768;
 end   
19'd153604: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=85;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1475;
 end   
19'd153605: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=37;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=669;
 end   
19'd153606: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=90;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=1580;
 end   
19'd153607: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=87;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=1539;
 end   
19'd153608: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=8;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=206;
 end   
19'd153609: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=85;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=1525;
 end   
19'd153610: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=42;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=804;
 end   
19'd153611: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=50;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=1715;
 end   
19'd153612: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=82;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=5691;
 end   
19'd153613: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=71;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=4318;
 end   
19'd153614: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=30;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=2975;
 end   
19'd153615: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=77;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=4519;
 end   
19'd153616: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=72;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=5180;
 end   
19'd153617: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=49;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=3989;
 end   
19'd153618: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=72;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=3806;
 end   
19'd153619: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=63;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=4675;
 end   
19'd153620: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=45;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=3054;
 end   
19'd153621: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd153763: begin  
rid<=1;
end
19'd153764: begin  
end
19'd153765: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd153766: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd153767: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd153768: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd153769: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd153770: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd153771: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd153772: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd153773: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd153774: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd153775: begin  
rid<=0;
end
19'd153901: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=84;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13964;
 end   
19'd153902: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=29;
   mapp<=64;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12098;
 end   
19'd153903: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=39;
   mapp<=50;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10870;
 end   
19'd153904: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=78;
   mapp<=99;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=8360;
 end   
19'd153905: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=49;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=8981;
 end   
19'd153906: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=23;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7934;
 end   
19'd153907: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=18;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd153908: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=52;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd153909: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=35;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd153910: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=11;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=28547;
 end   
19'd153911: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=73;
   mapp<=64;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=25063;
 end   
19'd153912: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=97;
   mapp<=38;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=26627;
 end   
19'd153913: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=89;
   mapp<=65;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=20961;
 end   
19'd153914: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=7;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=21207;
 end   
19'd153915: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=91;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=20794;
 end   
19'd153916: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=79;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd153917: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=48;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd153918: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=36;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd153919: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd154061: begin  
rid<=1;
end
19'd154062: begin  
end
19'd154063: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd154064: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd154065: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd154066: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd154067: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd154068: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd154069: begin  
rid<=0;
end
19'd154201: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=49;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12128;
 end   
19'd154202: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=58;
   mapp<=80;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8796;
 end   
19'd154203: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=17;
   mapp<=43;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8229;
 end   
19'd154204: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=35;
   mapp<=87;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7239;
 end   
19'd154205: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=8;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd154206: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd154207: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd154208: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd154209: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=82;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=24337;
 end   
19'd154210: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=25;
   mapp<=14;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=21488;
 end   
19'd154211: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=69;
   mapp<=20;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=23204;
 end   
19'd154212: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=2;
   mapp<=90;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=21648;
 end   
19'd154213: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=91;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd154214: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd154215: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd154216: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd154217: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd154359: begin  
rid<=1;
end
19'd154360: begin  
end
19'd154361: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd154362: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd154363: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd154364: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd154365: begin  
rid<=0;
end
19'd154501: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=37;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6680;
 end   
19'd154502: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=72;
   mapp<=15;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5940;
 end   
19'd154503: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=2;
   mapp<=43;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9400;
 end   
19'd154504: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=25;
   mapp<=77;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=10665;
 end   
19'd154505: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=85;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=11606;
 end   
19'd154506: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=83;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=9102;
 end   
19'd154507: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd154508: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd154509: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd154510: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=91;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=11018;
 end   
19'd154511: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=45;
   mapp<=25;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=14425;
 end   
19'd154512: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=66;
   mapp<=28;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=18953;
 end   
19'd154513: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=75;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=22671;
 end   
19'd154514: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=55;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=21954;
 end   
19'd154515: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=41;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=15878;
 end   
19'd154516: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd154517: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd154518: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd154519: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd154661: begin  
rid<=1;
end
19'd154662: begin  
end
19'd154663: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd154664: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd154665: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd154666: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd154667: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd154668: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd154669: begin  
rid<=0;
end
19'd154801: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=71;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7859;
 end   
19'd154802: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=69;
   mapp<=23;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7538;
 end   
19'd154803: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=57;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd154804: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=74;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd154805: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=12;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd154806: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd154807: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=68;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=21855;
 end   
19'd154808: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=96;
   mapp<=52;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=27640;
 end   
19'd154809: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=2;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd154810: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=98;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd154811: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=26;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd154812: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=87;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd154813: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd154955: begin  
rid<=1;
end
19'd154956: begin  
end
19'd154957: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd154958: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd154959: begin  
rid<=0;
end
19'd155101: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=91;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=20860;
 end   
19'd155102: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=94;
   mapp<=39;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=13627;
 end   
19'd155103: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=58;
   mapp<=18;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12848;
 end   
19'd155104: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=50;
   mapp<=17;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=15014;
 end   
19'd155105: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=69;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd155106: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=17;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd155107: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=23;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd155108: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=2;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd155109: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd155110: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=68;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd155111: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=33;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=47834;
 end   
19'd155112: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=52;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=39810;
 end   
19'd155113: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=17;
   mapp<=64;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=41127;
 end   
19'd155114: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=99;
   mapp<=39;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=47377;
 end   
19'd155115: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=89;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd155116: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=70;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd155117: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=85;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd155118: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=54;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd155119: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd155120: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=99;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd155121: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd155263: begin  
rid<=1;
end
19'd155264: begin  
end
19'd155265: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd155266: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd155267: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd155268: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd155269: begin  
rid<=0;
end
19'd155401: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=15;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4710;
 end   
19'd155402: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=45;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3205;
 end   
19'd155403: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=47;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3065;
 end   
19'd155404: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=52;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3330;
 end   
19'd155405: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=56;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1465;
 end   
19'd155406: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=13;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=605;
 end   
19'd155407: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd155408: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=40;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5226;
 end   
19'd155409: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=34;
   mapp<=14;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=6655;
 end   
19'd155410: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=85;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=7519;
 end   
19'd155411: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=31;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=5862;
 end   
19'd155412: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=38;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=3189;
 end   
19'd155413: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=6;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=2205;
 end   
19'd155414: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd155415: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd155557: begin  
rid<=1;
end
19'd155558: begin  
end
19'd155559: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd155560: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd155561: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd155562: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd155563: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd155564: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd155565: begin  
rid<=0;
end
19'd155701: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=89;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4450;
 end   
19'd155702: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=59;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5261;
 end   
19'd155703: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=64;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5716;
 end   
19'd155704: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=68;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6082;
 end   
19'd155705: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=12;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1108;
 end   
19'd155706: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=87;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7793;
 end   
19'd155707: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=46;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=4154;
 end   
19'd155708: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=74;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=6656;
 end   
19'd155709: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=98;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=8802;
 end   
19'd155710: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=6;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=4672;
 end   
19'd155711: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=20;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=5381;
 end   
19'd155712: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=95;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=6286;
 end   
19'd155713: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=14;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6166;
 end   
19'd155714: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=32;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=1300;
 end   
19'd155715: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=65;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=8183;
 end   
19'd155716: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=52;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=4466;
 end   
19'd155717: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=91;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=7202;
 end   
19'd155718: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=95;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=9372;
 end   
19'd155719: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd155861: begin  
rid<=1;
end
19'd155862: begin  
end
19'd155863: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd155864: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd155865: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd155866: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd155867: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd155868: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd155869: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd155870: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd155871: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd155872: begin  
rid<=0;
end
19'd156001: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=92;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6754;
 end   
19'd156002: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=52;
   mapp<=17;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9123;
 end   
19'd156003: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=19;
   mapp<=62;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6516;
 end   
19'd156004: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=99;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6629;
 end   
19'd156005: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd156006: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=8;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd156007: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=69;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14053;
 end   
19'd156008: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=57;
   mapp<=13;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=16218;
 end   
19'd156009: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=27;
   mapp<=18;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=11832;
 end   
19'd156010: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=96;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=17433;
 end   
19'd156011: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=94;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd156012: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=63;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd156013: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd156155: begin  
rid<=1;
end
19'd156156: begin  
end
19'd156157: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd156158: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd156159: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd156160: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd156161: begin  
rid<=0;
end
19'd156301: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=80;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8656;
 end   
19'd156302: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=72;
   mapp<=38;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10106;
 end   
19'd156303: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=98;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8292;
 end   
19'd156304: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=6;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=2670;
 end   
19'd156305: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=30;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5968;
 end   
19'd156306: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=49;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7714;
 end   
19'd156307: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=52;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=8324;
 end   
19'd156308: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=57;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=10678;
 end   
19'd156309: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd156310: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=79;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16720;
 end   
19'd156311: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=92;
   mapp<=43;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=19851;
 end   
19'd156312: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=69;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=16963;
 end   
19'd156313: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=35;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=13071;
 end   
19'd156314: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=83;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=14089;
 end   
19'd156315: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=17;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=13105;
 end   
19'd156316: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=44;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=12536;
 end   
19'd156317: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=8;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=14254;
 end   
19'd156318: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd156319: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd156461: begin  
rid<=1;
end
19'd156462: begin  
end
19'd156463: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd156464: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd156465: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd156466: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd156467: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd156468: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd156469: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd156470: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd156471: begin  
rid<=0;
end
19'd156601: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=61;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9585;
 end   
19'd156602: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=96;
   mapp<=3;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7515;
 end   
19'd156603: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=55;
   mapp<=21;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12472;
 end   
19'd156604: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=54;
   mapp<=25;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=12197;
 end   
19'd156605: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=27;
   mapp<=28;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=16201;
 end   
19'd156606: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=6;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd156607: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=34;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd156608: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd156609: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd156610: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd156611: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd156612: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=7;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=22049;
 end   
19'd156613: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=56;
   mapp<=19;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=23133;
 end   
19'd156614: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=47;
   mapp<=65;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=27788;
 end   
19'd156615: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=23;
   mapp<=83;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=26793;
 end   
19'd156616: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=20;
   mapp<=52;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=31913;
 end   
19'd156617: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=35;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd156618: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=47;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd156619: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd156620: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd156621: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd156622: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd156623: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd156765: begin  
rid<=1;
end
19'd156766: begin  
end
19'd156767: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd156768: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd156769: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd156770: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd156771: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd156772: begin  
rid<=0;
end
19'd156901: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=99;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16699;
 end   
19'd156902: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=80;
   mapp<=79;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=20956;
 end   
19'd156903: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=89;
   mapp<=1;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=16757;
 end   
19'd156904: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=9;
   mapp<=70;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=20518;
 end   
19'd156905: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=10;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd156906: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=34;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd156907: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=66;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd156908: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=62;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd156909: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=58;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd156910: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=22;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd156911: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=78;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd156912: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=10;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=32563;
 end   
19'd156913: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=97;
   mapp<=59;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=40556;
 end   
19'd156914: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=6;
   mapp<=37;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=35181;
 end   
19'd156915: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=47;
   mapp<=61;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=41834;
 end   
19'd156916: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=29;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd156917: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=63;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd156918: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=83;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd156919: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=4;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd156920: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=99;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd156921: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=85;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd156922: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=39;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd156923: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd157065: begin  
rid<=1;
end
19'd157066: begin  
end
19'd157067: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd157068: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd157069: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd157070: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd157071: begin  
rid<=0;
end
19'd157201: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=45;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4974;
 end   
19'd157202: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=66;
   mapp<=16;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6060;
 end   
19'd157203: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=21;
   mapp<=58;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9939;
 end   
19'd157204: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=55;
   mapp<=27;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4836;
 end   
19'd157205: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=17;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=11488;
 end   
19'd157206: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=94;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6567;
 end   
19'd157207: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=9;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=8329;
 end   
19'd157208: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd157209: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd157210: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd157211: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=29;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17891;
 end   
19'd157212: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=33;
   mapp<=39;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=23241;
 end   
19'd157213: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=54;
   mapp<=65;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=21808;
 end   
19'd157214: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=93;
   mapp<=87;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=13419;
 end   
19'd157215: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=99;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=17965;
 end   
19'd157216: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=19;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=11111;
 end   
19'd157217: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=19;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=18123;
 end   
19'd157218: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd157219: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd157220: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd157221: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd157363: begin  
rid<=1;
end
19'd157364: begin  
end
19'd157365: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd157366: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd157367: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd157368: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd157369: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd157370: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd157371: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd157372: begin  
rid<=0;
end
19'd157501: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=29;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10327;
 end   
19'd157502: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=79;
   mapp<=18;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9185;
 end   
19'd157503: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=75;
   mapp<=82;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6789;
 end   
19'd157504: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=29;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5333;
 end   
19'd157505: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=28;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6222;
 end   
19'd157506: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=30;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7005;
 end   
19'd157507: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=40;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=6851;
 end   
19'd157508: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=39;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=8912;
 end   
19'd157509: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd157510: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd157511: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=85;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17826;
 end   
19'd157512: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=72;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=22066;
 end   
19'd157513: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=88;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=19813;
 end   
19'd157514: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=77;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=18214;
 end   
19'd157515: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=88;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=16222;
 end   
19'd157516: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=35;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=11132;
 end   
19'd157517: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=16;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=10947;
 end   
19'd157518: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=38;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=17974;
 end   
19'd157519: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd157520: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd157521: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd157663: begin  
rid<=1;
end
19'd157664: begin  
end
19'd157665: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd157666: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd157667: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd157668: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd157669: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd157670: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd157671: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd157672: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd157673: begin  
rid<=0;
end
19'd157801: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=73;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10615;
 end   
19'd157802: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=70;
   mapp<=70;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6970;
 end   
19'd157803: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=16;
   mapp<=15;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5863;
 end   
19'd157804: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=50;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=9412;
 end   
19'd157805: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=78;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=8204;
 end   
19'd157806: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=17;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=8427;
 end   
19'd157807: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=80;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=12796;
 end   
19'd157808: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd157809: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd157810: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=75;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=24984;
 end   
19'd157811: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=35;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20356;
 end   
19'd157812: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=68;
   mapp<=93;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=18456;
 end   
19'd157813: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=42;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=20001;
 end   
19'd157814: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=61;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=19181;
 end   
19'd157815: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=78;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=16983;
 end   
19'd157816: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=54;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=20598;
 end   
19'd157817: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd157818: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd157819: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd157961: begin  
rid<=1;
end
19'd157962: begin  
end
19'd157963: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd157964: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd157965: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd157966: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd157967: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd157968: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd157969: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd157970: begin  
rid<=0;
end
19'd158101: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=23;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=21502;
 end   
19'd158102: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=57;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=25514;
 end   
19'd158103: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=72;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd158104: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=74;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd158105: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=58;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd158106: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=83;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd158107: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=4;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd158108: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=36;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=36149;
 end   
19'd158109: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=87;
   mapp<=16;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=44940;
 end   
19'd158110: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=30;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd158111: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=54;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd158112: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=35;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd158113: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=34;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd158114: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=78;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd158115: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd158257: begin  
rid<=1;
end
19'd158258: begin  
end
19'd158259: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd158260: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd158261: begin  
rid<=0;
end
19'd158401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=98;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16913;
 end   
19'd158402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=84;
   mapp<=12;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12996;
 end   
19'd158403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=16;
   mapp<=50;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=20396;
 end   
19'd158404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=26;
   mapp<=56;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=15710;
 end   
19'd158405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=64;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd158406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=7;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd158407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=51;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd158408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=10;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd158409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd158410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd158411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd158412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=39;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=38656;
 end   
19'd158413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=59;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=36305;
 end   
19'd158414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=67;
   mapp<=51;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=43432;
 end   
19'd158415: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=40;
   mapp<=20;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=37406;
 end   
19'd158416: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=25;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd158417: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=78;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd158418: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=28;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd158419: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=7;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd158420: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd158421: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd158422: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd158423: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd158565: begin  
rid<=1;
end
19'd158566: begin  
end
19'd158567: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd158568: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd158569: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd158570: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd158571: begin  
rid<=0;
end
19'd158701: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=81;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12584;
 end   
19'd158702: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=21;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=13996;
 end   
19'd158703: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=89;
   mapp<=58;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10988;
 end   
19'd158704: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=57;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=11985;
 end   
19'd158705: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=57;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=8064;
 end   
19'd158706: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=69;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6457;
 end   
19'd158707: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd158708: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd158709: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=47;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=15367;
 end   
19'd158710: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=14;
   mapp<=73;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=19061;
 end   
19'd158711: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=13;
   mapp<=74;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15175;
 end   
19'd158712: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=46;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=14529;
 end   
19'd158713: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=5;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=9519;
 end   
19'd158714: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=24;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=8576;
 end   
19'd158715: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd158716: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd158717: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd158859: begin  
rid<=1;
end
19'd158860: begin  
end
19'd158861: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd158862: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd158863: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd158864: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd158865: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd158866: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd158867: begin  
rid<=0;
end
19'd159001: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=9;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=24625;
 end   
19'd159002: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=13;
   mapp<=99;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=25371;
 end   
19'd159003: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=52;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd159004: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=93;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd159005: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=75;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd159006: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=56;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd159007: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=72;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd159008: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=26;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd159009: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=31;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=53528;
 end   
19'd159010: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=99;
   mapp<=86;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=58298;
 end   
19'd159011: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=96;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd159012: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=53;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd159013: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=70;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd159014: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=22;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd159015: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=75;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd159016: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=55;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd159017: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd159159: begin  
rid<=1;
end
19'd159160: begin  
end
19'd159161: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd159162: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd159163: begin  
rid<=0;
end
19'd159301: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=10;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=19824;
 end   
19'd159302: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=29;
   mapp<=66;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=17016;
 end   
19'd159303: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=34;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd159304: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=35;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd159305: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=70;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd159306: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=86;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd159307: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=5;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd159308: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=31;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd159309: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=23;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd159310: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=20;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd159311: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd159312: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=13;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=49104;
 end   
19'd159313: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=68;
   mapp<=82;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=40490;
 end   
19'd159314: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=12;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd159315: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=8;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd159316: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=46;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd159317: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=47;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd159318: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd159319: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=94;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd159320: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=96;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd159321: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=43;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd159322: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd159323: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd159465: begin  
rid<=1;
end
19'd159466: begin  
end
19'd159467: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd159468: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd159469: begin  
rid<=0;
end
19'd159601: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=94;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14669;
 end   
19'd159602: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=98;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd159603: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=25;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd159604: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=89;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd159605: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=55;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd159606: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=55;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd159607: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=42;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=39765;
 end   
19'd159608: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=88;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd159609: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=98;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd159610: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=94;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd159611: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=60;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd159612: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=98;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd159613: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd159755: begin  
rid<=1;
end
19'd159756: begin  
end
19'd159757: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd159758: begin  
rid<=0;
end
19'd159901: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=46;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7186;
 end   
19'd159902: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=97;
   mapp<=47;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10136;
 end   
19'd159903: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=15;
   mapp<=77;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7543;
 end   
19'd159904: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=33;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6742;
 end   
19'd159905: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=52;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3882;
 end   
19'd159906: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd159907: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd159908: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=40;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=11541;
 end   
19'd159909: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=52;
   mapp<=54;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=13497;
 end   
19'd159910: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=17;
   mapp<=11;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=11233;
 end   
19'd159911: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=37;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=12856;
 end   
19'd159912: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=78;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=9025;
 end   
19'd159913: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd159914: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd159915: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd160057: begin  
rid<=1;
end
19'd160058: begin  
end
19'd160059: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd160060: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd160061: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd160062: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd160063: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd160064: begin  
rid<=0;
end
19'd160201: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=23;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10017;
 end   
19'd160202: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=7;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8282;
 end   
19'd160203: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=48;
   mapp<=68;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=14006;
 end   
19'd160204: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=14;
   mapp<=37;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=10062;
 end   
19'd160205: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=71;
   mapp<=77;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=10781;
 end   
19'd160206: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=18;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=10327;
 end   
19'd160207: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=90;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=10399;
 end   
19'd160208: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=7;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd160209: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=29;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd160210: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=32;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd160211: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=72;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd160212: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=7;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=30699;
 end   
19'd160213: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=85;
   mapp<=87;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=29291;
 end   
19'd160214: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=84;
   mapp<=95;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=33556;
 end   
19'd160215: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=27;
   mapp<=87;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=29414;
 end   
19'd160216: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=44;
   mapp<=58;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=30176;
 end   
19'd160217: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=41;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=30168;
 end   
19'd160218: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=79;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=30400;
 end   
19'd160219: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=55;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd160220: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=17;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd160221: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=67;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd160222: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=55;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd160223: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd160365: begin  
rid<=1;
end
19'd160366: begin  
end
19'd160367: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd160368: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd160369: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd160370: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd160371: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd160372: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd160373: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd160374: begin  
rid<=0;
end
19'd160501: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=13;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=17860;
 end   
19'd160502: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=2;
   mapp<=69;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15057;
 end   
19'd160503: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=51;
   mapp<=60;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=14193;
 end   
19'd160504: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=75;
   mapp<=25;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=19033;
 end   
19'd160505: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=54;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd160506: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=67;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd160507: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=89;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd160508: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd160509: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd160510: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd160511: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=98;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=42895;
 end   
19'd160512: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=3;
   mapp<=61;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=41113;
 end   
19'd160513: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=41;
   mapp<=98;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=47055;
 end   
19'd160514: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=87;
   mapp<=48;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=48217;
 end   
19'd160515: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=86;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd160516: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=94;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd160517: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=88;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd160518: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd160519: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd160520: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd160521: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd160663: begin  
rid<=1;
end
19'd160664: begin  
end
19'd160665: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd160666: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd160667: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd160668: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd160669: begin  
rid<=0;
end
19'd160801: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=93;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8463;
 end   
19'd160802: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=90;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8200;
 end   
19'd160803: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=89;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8119;
 end   
19'd160804: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=92;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=8402;
 end   
19'd160805: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=15;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1405;
 end   
19'd160806: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=65;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=5965;
 end   
19'd160807: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=81;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=15024;
 end   
19'd160808: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=89;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=15409;
 end   
19'd160809: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=36;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=11035;
 end   
19'd160810: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=2;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=8564;
 end   
19'd160811: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=27;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=3592;
 end   
19'd160812: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=87;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=13012;
 end   
19'd160813: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd160955: begin  
rid<=1;
end
19'd160956: begin  
end
19'd160957: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd160958: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd160959: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd160960: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd160961: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd160962: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd160963: begin  
rid<=0;
end
19'd161101: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=53;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5471;
 end   
19'd161102: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=85;
   mapp<=7;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8418;
 end   
19'd161103: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=84;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7853;
 end   
19'd161104: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=15;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=2103;
 end   
19'd161105: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=99;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd161106: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=32;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=9077;
 end   
19'd161107: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=47;
   mapp<=74;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=10012;
 end   
19'd161108: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=19;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=10149;
 end   
19'd161109: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=30;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=9549;
 end   
19'd161110: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=99;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd161111: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd161253: begin  
rid<=1;
end
19'd161254: begin  
end
19'd161255: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd161256: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd161257: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd161258: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd161259: begin  
rid<=0;
end
19'd161401: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=62;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6091;
 end   
19'd161402: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=71;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd161403: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=61;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=9766;
 end   
19'd161404: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=49;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd161405: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd161547: begin  
rid<=1;
end
19'd161548: begin  
end
19'd161549: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd161550: begin  
rid<=0;
end
19'd161701: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=13;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=52;
 end   
19'd161702: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=12;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=166;
 end   
19'd161703: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=42;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=566;
 end   
19'd161704: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=24;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=342;
 end   
19'd161705: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=19;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=287;
 end   
19'd161706: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=13;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=219;
 end   
19'd161707: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=42;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=606;
 end   
19'd161708: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=54;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=772;
 end   
19'd161709: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=65;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=925;
 end   
19'd161710: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=96;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=1338;
 end   
19'd161711: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=73;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=2169;
 end   
19'd161712: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=13;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=1115;
 end   
19'd161713: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=32;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=2902;
 end   
19'd161714: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=12;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=1218;
 end   
19'd161715: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=90;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=6857;
 end   
19'd161716: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=97;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=7300;
 end   
19'd161717: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=78;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=6300;
 end   
19'd161718: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=1;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=845;
 end   
19'd161719: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=4;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=1217;
 end   
19'd161720: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=8;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=1922;
 end   
19'd161721: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd161863: begin  
rid<=1;
end
19'd161864: begin  
end
19'd161865: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd161866: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd161867: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd161868: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd161869: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd161870: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd161871: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd161872: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd161873: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd161874: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd161875: begin  
rid<=0;
end
19'd162001: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=14;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6760;
 end   
19'd162002: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=55;
   mapp<=53;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11527;
 end   
19'd162003: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=5;
   mapp<=92;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7318;
 end   
19'd162004: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=75;
   mapp<=33;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=8717;
 end   
19'd162005: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=74;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4891;
 end   
19'd162006: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd162007: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd162008: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd162009: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=71;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16390;
 end   
19'd162010: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=2;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18910;
 end   
19'd162011: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=14;
   mapp<=77;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=16745;
 end   
19'd162012: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=58;
   mapp<=54;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=19035;
 end   
19'd162013: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=10;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=10495;
 end   
19'd162014: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd162015: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd162016: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd162017: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd162159: begin  
rid<=1;
end
19'd162160: begin  
end
19'd162161: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd162162: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd162163: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd162164: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd162165: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd162166: begin  
rid<=0;
end
19'd162301: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=41;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7398;
 end   
19'd162302: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=60;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11114;
 end   
19'd162303: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=24;
   mapp<=38;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12648;
 end   
19'd162304: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=20;
   mapp<=96;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=10476;
 end   
19'd162305: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=86;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=15062;
 end   
19'd162306: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=81;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=5748;
 end   
19'd162307: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=11;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=10038;
 end   
19'd162308: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=86;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=3222;
 end   
19'd162309: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd162310: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd162311: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=5;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd162312: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=25;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16070;
 end   
19'd162313: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=45;
   mapp<=4;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18896;
 end   
19'd162314: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=65;
   mapp<=78;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=19934;
 end   
19'd162315: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=38;
   mapp<=44;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=14608;
 end   
19'd162316: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=32;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=19504;
 end   
19'd162317: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=2;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=8836;
 end   
19'd162318: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=27;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=21050;
 end   
19'd162319: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=2;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=15332;
 end   
19'd162320: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=61;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd162321: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=99;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd162322: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=91;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd162323: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd162465: begin  
rid<=1;
end
19'd162466: begin  
end
19'd162467: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd162468: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd162469: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd162470: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd162471: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd162472: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd162473: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd162474: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd162475: begin  
rid<=0;
end
19'd162601: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=42;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2745;
 end   
19'd162602: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=15;
   mapp<=3;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3214;
 end   
19'd162603: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=36;
   mapp<=54;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6797;
 end   
19'd162604: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd162605: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd162606: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=40;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8287;
 end   
19'd162607: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=6;
   mapp<=26;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12399;
 end   
19'd162608: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=99;
   mapp<=54;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=18935;
 end   
19'd162609: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd162610: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd162611: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd162753: begin  
rid<=1;
end
19'd162754: begin  
end
19'd162755: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd162756: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd162757: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd162758: begin  
rid<=0;
end
19'd162901: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=83;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5662;
 end   
19'd162902: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=29;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd162903: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=9;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7435;
 end   
19'd162904: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=20;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd162905: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd163047: begin  
rid<=1;
end
19'd163048: begin  
end
19'd163049: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd163050: begin  
rid<=0;
end
19'd163201: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=99;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1881;
 end   
19'd163202: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=68;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1302;
 end   
19'd163203: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=56;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1084;
 end   
19'd163204: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=23;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=467;
 end   
19'd163205: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=30;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=610;
 end   
19'd163206: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=18;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=392;
 end   
19'd163207: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=17;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=383;
 end   
19'd163208: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=2;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=108;
 end   
19'd163209: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=34;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=4499;
 end   
19'd163210: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=68;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=6538;
 end   
19'd163211: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=23;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=2855;
 end   
19'd163212: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=41;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=3624;
 end   
19'd163213: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=81;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=6847;
 end   
19'd163214: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=78;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=6398;
 end   
19'd163215: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=82;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=6697;
 end   
19'd163216: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=7;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=647;
 end   
19'd163217: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd163359: begin  
rid<=1;
end
19'd163360: begin  
end
19'd163361: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd163362: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd163363: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd163364: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd163365: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd163366: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd163367: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd163368: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd163369: begin  
rid<=0;
end
19'd163501: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=8;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=18128;
 end   
19'd163502: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=26;
   mapp<=33;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=17525;
 end   
19'd163503: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=39;
   mapp<=21;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=16139;
 end   
19'd163504: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=76;
   mapp<=80;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=20981;
 end   
19'd163505: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=87;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd163506: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd163507: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=57;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd163508: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=70;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd163509: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=20;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd163510: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=51;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd163511: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=24;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd163512: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=86;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=42221;
 end   
19'd163513: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=17;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=34056;
 end   
19'd163514: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=1;
   mapp<=80;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=32347;
 end   
19'd163515: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=46;
   mapp<=32;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=46515;
 end   
19'd163516: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=68;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd163517: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=76;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd163518: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=17;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd163519: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=56;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd163520: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=1;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd163521: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd163522: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=84;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd163523: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd163665: begin  
rid<=1;
end
19'd163666: begin  
end
19'd163667: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd163668: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd163669: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd163670: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd163671: begin  
rid<=0;
end
19'd163801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=56;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6465;
 end   
19'd163802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=6;
   mapp<=61;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4833;
 end   
19'd163803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=17;
   mapp<=13;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8048;
 end   
19'd163804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=32;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd163805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=5;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd163806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=33;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd163807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd163808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=78;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd163809: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=34;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=20588;
 end   
19'd163810: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=1;
   mapp<=30;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=17844;
 end   
19'd163811: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=73;
   mapp<=90;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=19635;
 end   
19'd163812: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=33;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd163813: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=36;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd163814: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=12;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd163815: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=53;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd163816: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=5;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd163817: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd163959: begin  
rid<=1;
end
19'd163960: begin  
end
19'd163961: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd163962: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd163963: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd163964: begin  
rid<=0;
end
19'd164101: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=22;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7656;
 end   
19'd164102: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=48;
   mapp<=47;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5761;
 end   
19'd164103: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=3;
   mapp<=35;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11187;
 end   
19'd164104: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=96;
   mapp<=45;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=16252;
 end   
19'd164105: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=1;
   mapp<=95;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=10541;
 end   
19'd164106: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=3;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=9944;
 end   
19'd164107: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=67;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd164108: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=97;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd164109: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd164110: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd164111: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=32;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=22102;
 end   
19'd164112: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=75;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=21622;
 end   
19'd164113: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=67;
   mapp<=0;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=23143;
 end   
19'd164114: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=35;
   mapp<=95;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=29539;
 end   
19'd164115: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=49;
   mapp<=50;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=17178;
 end   
19'd164116: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=20;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=22314;
 end   
19'd164117: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=65;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd164118: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=14;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd164119: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=17;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd164120: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=73;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd164121: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd164263: begin  
rid<=1;
end
19'd164264: begin  
end
19'd164265: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd164266: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd164267: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd164268: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd164269: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd164270: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd164271: begin  
rid<=0;
end
19'd164401: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=36;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4104;
 end   
19'd164402: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=58;
   mapp<=54;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6868;
 end   
19'd164403: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=98;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6608;
 end   
19'd164404: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=73;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4215;
 end   
19'd164405: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=41;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2389;
 end   
19'd164406: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=23;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=2129;
 end   
19'd164407: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=27;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=5919;
 end   
19'd164408: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=95;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=3121;
 end   
19'd164409: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=9;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd164410: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=23;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=10981;
 end   
19'd164411: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=69;
   mapp<=71;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=17346;
 end   
19'd164412: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=64;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=16017;
 end   
19'd164413: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=55;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=11359;
 end   
19'd164414: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=34;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=12058;
 end   
19'd164415: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=95;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=14062;
 end   
19'd164416: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=53;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=15731;
 end   
19'd164417: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=74;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=10905;
 end   
19'd164418: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=20;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd164419: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd164561: begin  
rid<=1;
end
19'd164562: begin  
end
19'd164563: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd164564: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd164565: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd164566: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd164567: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd164568: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd164569: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd164570: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd164571: begin  
rid<=0;
end
19'd164701: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=24;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5155;
 end   
19'd164702: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=76;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd164703: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=39;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd164704: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=71;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd164705: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=30;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12017;
 end   
19'd164706: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=21;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd164707: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=10;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd164708: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=85;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd164709: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd164851: begin  
rid<=1;
end
19'd164852: begin  
end
19'd164853: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd164854: begin  
rid<=0;
end
19'd165001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=2;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11482;
 end   
19'd165002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=87;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4255;
 end   
19'd165003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=30;
   mapp<=5;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10844;
 end   
19'd165004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=47;
   mapp<=87;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6447;
 end   
19'd165005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=22;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=10010;
 end   
19'd165006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=55;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=10317;
 end   
19'd165007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=57;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=11312;
 end   
19'd165008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=73;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=10152;
 end   
19'd165009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd165010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd165011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd165012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=43;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=15296;
 end   
19'd165013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=79;
   mapp<=28;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=11447;
 end   
19'd165014: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=6;
   mapp<=51;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=14593;
 end   
19'd165015: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=25;
   mapp<=14;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=13149;
 end   
19'd165016: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=75;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=15502;
 end   
19'd165017: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=12954;
 end   
19'd165018: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=7;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=19641;
 end   
19'd165019: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=89;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=19202;
 end   
19'd165020: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd165021: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd165022: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd165023: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd165165: begin  
rid<=1;
end
19'd165166: begin  
end
19'd165167: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd165168: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd165169: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd165170: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd165171: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd165172: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd165173: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd165174: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd165175: begin  
rid<=0;
end
19'd165301: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=50;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5705;
 end   
19'd165302: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=51;
   mapp<=20;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5756;
 end   
19'd165303: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=29;
   mapp<=9;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5400;
 end   
19'd165304: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=60;
   mapp<=19;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7784;
 end   
19'd165305: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=1;
   mapp<=34;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4714;
 end   
19'd165306: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=38;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7989;
 end   
19'd165307: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=46;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd165308: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=77;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd165309: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=58;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd165310: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=81;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd165311: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=59;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=11687;
 end   
19'd165312: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=15;
   mapp<=37;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=9414;
 end   
19'd165313: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=59;
   mapp<=7;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=12105;
 end   
19'd165314: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=55;
   mapp<=3;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=15782;
 end   
19'd165315: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=89;
   mapp<=22;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=10826;
 end   
19'd165316: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=4;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=12849;
 end   
19'd165317: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=52;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd165318: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=83;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd165319: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=45;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd165320: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=92;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd165321: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd165463: begin  
rid<=1;
end
19'd165464: begin  
end
19'd165465: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd165466: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd165467: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd165468: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd165469: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd165470: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd165471: begin  
rid<=0;
end
19'd165601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=21;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6156;
 end   
19'd165602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=78;
   mapp<=20;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9201;
 end   
19'd165603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=7;
   mapp<=64;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5393;
 end   
19'd165604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=31;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd165605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=35;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd165606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd165607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd165608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=92;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=21225;
 end   
19'd165609: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=83;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=25183;
 end   
19'd165610: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=31;
   mapp<=89;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=22045;
 end   
19'd165611: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=22;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd165612: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=48;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd165613: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd165614: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd165615: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd165757: begin  
rid<=1;
end
19'd165758: begin  
end
19'd165759: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd165760: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd165761: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd165762: begin  
rid<=0;
end
19'd165901: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=56;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=22434;
 end   
19'd165902: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=36;
   mapp<=28;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=24200;
 end   
19'd165903: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=97;
   mapp<=68;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=23039;
 end   
19'd165904: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=77;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd165905: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=63;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd165906: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=38;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd165907: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=37;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd165908: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=10;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd165909: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd165910: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd165911: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=24;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=42203;
 end   
19'd165912: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=54;
   mapp<=64;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=49428;
 end   
19'd165913: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=8;
   mapp<=78;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=46015;
 end   
19'd165914: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd165915: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=86;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd165916: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=67;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd165917: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=78;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd165918: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=50;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd165919: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd165920: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd165921: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd166063: begin  
rid<=1;
end
19'd166064: begin  
end
19'd166065: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd166066: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd166067: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd166068: begin  
rid<=0;
end
19'd166201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=87;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8436;
 end   
19'd166202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=19;
   mapp<=9;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=850;
 end   
19'd166203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd166204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=70;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14090;
 end   
19'd166205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=22;
   mapp<=82;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8768;
 end   
19'd166206: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd166207: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd166349: begin  
rid<=1;
end
19'd166350: begin  
end
19'd166351: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd166352: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd166353: begin  
rid<=0;
end
19'd166501: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=51;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10383;
 end   
19'd166502: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=2;
   mapp<=39;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8127;
 end   
19'd166503: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=59;
   mapp<=42;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9973;
 end   
19'd166504: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=20;
   mapp<=42;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=8883;
 end   
19'd166505: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=51;
   mapp<=80;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=11487;
 end   
19'd166506: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd166507: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=28;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd166508: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=39;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd166509: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=55;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd166510: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=58;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14429;
 end   
19'd166511: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=3;
   mapp<=39;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=16343;
 end   
19'd166512: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=10;
   mapp<=76;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=17102;
 end   
19'd166513: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=66;
   mapp<=19;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=18613;
 end   
19'd166514: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=5;
   mapp<=35;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=22267;
 end   
19'd166515: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=75;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd166516: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd166517: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=15;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd166518: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=60;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd166519: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd166661: begin  
rid<=1;
end
19'd166662: begin  
end
19'd166663: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd166664: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd166665: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd166666: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd166667: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd166668: begin  
rid<=0;
end
19'd166801: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=55;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14000;
 end   
19'd166802: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=15;
   mapp<=57;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15236;
 end   
19'd166803: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=95;
   mapp<=69;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=16017;
 end   
19'd166804: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=35;
   mapp<=83;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=11684;
 end   
19'd166805: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=77;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=9279;
 end   
19'd166806: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=28;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=4310;
 end   
19'd166807: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=36;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd166808: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd166809: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=4;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd166810: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=13;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16557;
 end   
19'd166811: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=52;
   mapp<=1;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=21660;
 end   
19'd166812: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=37;
   mapp<=28;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=22275;
 end   
19'd166813: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=26;
   mapp<=7;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=16669;
 end   
19'd166814: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=73;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=17561;
 end   
19'd166815: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=75;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=11902;
 end   
19'd166816: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd166817: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=4;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd166818: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=3;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd166819: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd166961: begin  
rid<=1;
end
19'd166962: begin  
end
19'd166963: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd166964: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd166965: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd166966: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd166967: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd166968: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd166969: begin  
rid<=0;
end
19'd167101: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=21;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3971;
 end   
19'd167102: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=83;
   mapp<=11;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4751;
 end   
19'd167103: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=97;
   mapp<=22;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5399;
 end   
19'd167104: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=1;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=2516;
 end   
19'd167105: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=50;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd167106: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=86;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd167107: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=64;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12944;
 end   
19'd167108: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=96;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=11510;
 end   
19'd167109: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=53;
   mapp<=89;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=14394;
 end   
19'd167110: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=40;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=12090;
 end   
19'd167111: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=77;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd167112: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=71;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd167113: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd167255: begin  
rid<=1;
end
19'd167256: begin  
end
19'd167257: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd167258: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd167259: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd167260: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd167261: begin  
rid<=0;
end
19'd167401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=50;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9661;
 end   
19'd167402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=76;
   mapp<=45;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15704;
 end   
19'd167403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=80;
   mapp<=28;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11184;
 end   
19'd167404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=21;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd167405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=5;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd167406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=42;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd167407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd167408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd167409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=14;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=22613;
 end   
19'd167410: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=67;
   mapp<=52;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=33332;
 end   
19'd167411: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=94;
   mapp<=4;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=27632;
 end   
19'd167412: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=92;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd167413: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=44;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd167414: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=80;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd167415: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd167416: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd167417: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd167559: begin  
rid<=1;
end
19'd167560: begin  
end
19'd167561: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd167562: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd167563: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd167564: begin  
rid<=0;
end
19'd167701: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=40;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11041;
 end   
19'd167702: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=24;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10329;
 end   
19'd167703: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=63;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd167704: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=34;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd167705: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=53;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd167706: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=5;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd167707: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd167708: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=93;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=31523;
 end   
19'd167709: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=45;
   mapp<=81;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=31256;
 end   
19'd167710: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=53;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd167711: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=86;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd167712: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=22;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd167713: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=87;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd167714: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd167715: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd167857: begin  
rid<=1;
end
19'd167858: begin  
end
19'd167859: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd167860: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd167861: begin  
rid<=0;
end
19'd168001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=92;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4693;
 end   
19'd168002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=38;
   mapp<=49;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3105;
 end   
19'd168003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=29;
   mapp<=60;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2443;
 end   
19'd168004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=10;
   mapp<=28;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4030;
 end   
19'd168005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=5;
   mapp<=15;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5025;
 end   
19'd168006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=42;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6109;
 end   
19'd168007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=15;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=6916;
 end   
19'd168008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=49;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd168009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=41;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd168010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=60;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd168011: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=13;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd168012: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=94;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=13883;
 end   
19'd168013: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=81;
   mapp<=3;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=16485;
 end   
19'd168014: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=38;
   mapp<=81;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=10186;
 end   
19'd168015: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=75;
   mapp<=1;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=13734;
 end   
19'd168016: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=26;
   mapp<=71;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=13084;
 end   
19'd168017: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=53;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=12734;
 end   
19'd168018: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=53;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=17417;
 end   
19'd168019: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=30;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd168020: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=35;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd168021: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=25;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd168022: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=75;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd168023: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd168165: begin  
rid<=1;
end
19'd168166: begin  
end
19'd168167: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd168168: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd168169: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd168170: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd168171: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd168172: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd168173: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd168174: begin  
rid<=0;
end
19'd168301: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=4;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2510;
 end   
19'd168302: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=26;
   mapp<=89;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2264;
 end   
19'd168303: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd168304: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=88;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5766;
 end   
19'd168305: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=33;
   mapp<=64;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8556;
 end   
19'd168306: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd168307: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd168449: begin  
rid<=1;
end
19'd168450: begin  
end
19'd168451: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd168452: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd168453: begin  
rid<=0;
end
19'd168601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=48;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11768;
 end   
19'd168602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=56;
   mapp<=61;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9722;
 end   
19'd168603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=59;
   mapp<=33;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6729;
 end   
19'd168604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=87;
   mapp<=35;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=12649;
 end   
19'd168605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd168606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd168607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd168608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=28;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17189;
 end   
19'd168609: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=18;
   mapp<=27;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=14336;
 end   
19'd168610: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=34;
   mapp<=7;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=11928;
 end   
19'd168611: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=35;
   mapp<=83;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=20406;
 end   
19'd168612: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd168613: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd168614: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd168615: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd168757: begin  
rid<=1;
end
19'd168758: begin  
end
19'd168759: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd168760: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd168761: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd168762: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd168763: begin  
rid<=0;
end
19'd168901: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=28;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=420;
 end   
19'd168902: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=23;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=654;
 end   
19'd168903: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=85;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2400;
 end   
19'd168904: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=77;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=2186;
 end   
19'd168905: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=40;
 end   
19'd168906: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=25;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=750;
 end   
19'd168907: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=56;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=1628;
 end   
19'd168908: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=36;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=1078;
 end   
19'd168909: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=38;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=1144;
 end   
19'd168910: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=61;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=1518;
 end   
19'd168911: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=19;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=1813;
 end   
19'd168912: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=49;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=5389;
 end   
19'd168913: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=3;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=2369;
 end   
19'd168914: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=46;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=2846;
 end   
19'd168915: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=52;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=3922;
 end   
19'd168916: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=9;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=2177;
 end   
19'd168917: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=11;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=1749;
 end   
19'd168918: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=59;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=4743;
 end   
19'd168919: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd169061: begin  
rid<=1;
end
19'd169062: begin  
end
19'd169063: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd169064: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd169065: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd169066: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd169067: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd169068: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd169069: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd169070: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd169071: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd169072: begin  
rid<=0;
end
19'd169201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=24;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7766;
 end   
19'd169202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=14;
   mapp<=76;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11913;
 end   
19'd169203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=91;
   mapp<=60;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8903;
 end   
19'd169204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=70;
   mapp<=15;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5405;
 end   
19'd169205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=45;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5014;
 end   
19'd169206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=9;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6524;
 end   
19'd169207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=57;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd169208: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd169209: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=2;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd169210: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=55;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17219;
 end   
19'd169211: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=77;
   mapp<=18;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=19398;
 end   
19'd169212: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=67;
   mapp<=60;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=17054;
 end   
19'd169213: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=23;
   mapp<=54;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=15740;
 end   
19'd169214: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=18;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=16504;
 end   
19'd169215: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=60;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=16706;
 end   
19'd169216: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=97;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd169217: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=68;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd169218: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=24;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd169219: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd169361: begin  
rid<=1;
end
19'd169362: begin  
end
19'd169363: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd169364: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd169365: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd169366: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd169367: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd169368: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd169369: begin  
rid<=0;
end
19'd169501: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=31;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12859;
 end   
19'd169502: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=75;
   mapp<=96;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11864;
 end   
19'd169503: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=41;
   mapp<=73;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11501;
 end   
19'd169504: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=83;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=8119;
 end   
19'd169505: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=73;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3526;
 end   
19'd169506: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=1;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=4682;
 end   
19'd169507: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=28;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=8496;
 end   
19'd169508: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd169509: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd169510: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=16;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=19250;
 end   
19'd169511: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=39;
   mapp<=73;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18666;
 end   
19'd169512: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=90;
   mapp<=36;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=17330;
 end   
19'd169513: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=47;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=16113;
 end   
19'd169514: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=38;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=12930;
 end   
19'd169515: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=64;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=12846;
 end   
19'd169516: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=70;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=19897;
 end   
19'd169517: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd169518: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd169519: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd169661: begin  
rid<=1;
end
19'd169662: begin  
end
19'd169663: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd169664: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd169665: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd169666: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd169667: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd169668: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd169669: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd169670: begin  
rid<=0;
end
19'd169801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=21;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=17661;
 end   
19'd169802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=65;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=22433;
 end   
19'd169803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=33;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd169804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=92;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd169805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=63;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd169806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=13;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd169807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=98;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd169808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=90;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=32610;
 end   
19'd169809: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=75;
   mapp<=16;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=33594;
 end   
19'd169810: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=85;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd169811: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=77;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd169812: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=19;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd169813: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=3;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd169814: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=45;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd169815: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd169957: begin  
rid<=1;
end
19'd169958: begin  
end
19'd169959: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd169960: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd169961: begin  
rid<=0;
end
19'd170101: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=7;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4154;
 end   
19'd170102: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=38;
   mapp<=96;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5264;
 end   
19'd170103: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=37;
   mapp<=2;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9008;
 end   
19'd170104: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=76;
   mapp<=2;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4850;
 end   
19'd170105: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=15;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd170106: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=91;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd170107: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=79;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd170108: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=92;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7603;
 end   
19'd170109: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=55;
   mapp<=6;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=11830;
 end   
19'd170110: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=31;
   mapp<=65;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=11793;
 end   
19'd170111: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=88;
   mapp<=0;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=10500;
 end   
19'd170112: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=29;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd170113: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=68;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd170114: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=48;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd170115: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd170257: begin  
rid<=1;
end
19'd170258: begin  
end
19'd170259: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd170260: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd170261: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd170262: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd170263: begin  
rid<=0;
end
19'd170401: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=99;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12141;
 end   
19'd170402: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=36;
   mapp<=65;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4549;
 end   
19'd170403: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=15;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6185;
 end   
19'd170404: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=72;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=8068;
 end   
19'd170405: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=14;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd170406: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=78;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=19325;
 end   
19'd170407: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=80;
   mapp<=4;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=11689;
 end   
19'd170408: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=25;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=8537;
 end   
19'd170409: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=38;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=11704;
 end   
19'd170410: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=73;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd170411: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd170553: begin  
rid<=1;
end
19'd170554: begin  
end
19'd170555: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd170556: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd170557: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd170558: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd170559: begin  
rid<=0;
end
19'd170701: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=91;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1274;
 end   
19'd170702: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=25;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2285;
 end   
19'd170703: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=4;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=384;
 end   
19'd170704: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=1;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=121;
 end   
19'd170705: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=73;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6683;
 end   
19'd170706: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=63;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=5783;
 end   
19'd170707: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=58;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=5338;
 end   
19'd170708: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=50;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=4620;
 end   
19'd170709: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=59;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=3634;
 end   
19'd170710: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=17;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=3288;
 end   
19'd170711: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=29;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=2095;
 end   
19'd170712: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=28;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=1773;
 end   
19'd170713: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=81;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=11462;
 end   
19'd170714: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=53;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=8910;
 end   
19'd170715: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=84;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=10294;
 end   
19'd170716: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=4;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=4856;
 end   
19'd170717: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd170859: begin  
rid<=1;
end
19'd170860: begin  
end
19'd170861: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd170862: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd170863: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd170864: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd170865: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd170866: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd170867: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd170868: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd170869: begin  
rid<=0;
end
19'd171001: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=6;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1763;
 end   
19'd171002: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=55;
   mapp<=29;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3116;
 end   
19'd171003: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=54;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3011;
 end   
19'd171004: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=51;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3981;
 end   
19'd171005: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=87;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4709;
 end   
19'd171006: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=77;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=5019;
 end   
19'd171007: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=97;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=4429;
 end   
19'd171008: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=57;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=2710;
 end   
19'd171009: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=36;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=2248;
 end   
19'd171010: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=40;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=1964;
 end   
19'd171011: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=26;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd171012: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=4;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=2051;
 end   
19'd171013: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=26;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=4988;
 end   
19'd171014: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=25;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=4811;
 end   
19'd171015: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=53;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=7797;
 end   
19'd171016: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=64;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=9317;
 end   
19'd171017: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=98;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=12075;
 end   
19'd171018: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=16;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=5581;
 end   
19'd171019: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=63;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=7246;
 end   
19'd171020: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=94;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=9016;
 end   
19'd171021: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=19;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=3332;
 end   
19'd171022: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=42;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd171023: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd171165: begin  
rid<=1;
end
19'd171166: begin  
end
19'd171167: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd171168: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd171169: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd171170: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd171171: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd171172: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd171173: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd171174: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd171175: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd171176: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd171177: begin  
rid<=0;
end
19'd171301: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=95;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=20906;
 end   
19'd171302: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=33;
   mapp<=30;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=23221;
 end   
19'd171303: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=80;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd171304: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=18;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd171305: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=13;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd171306: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=70;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd171307: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=36;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd171308: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=73;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd171309: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=36;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd171310: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd171311: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=48;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=30774;
 end   
19'd171312: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=81;
   mapp<=17;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=40281;
 end   
19'd171313: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=9;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd171314: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=53;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd171315: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=31;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd171316: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=19;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd171317: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=52;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd171318: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=95;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd171319: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=3;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd171320: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd171321: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd171463: begin  
rid<=1;
end
19'd171464: begin  
end
19'd171465: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd171466: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd171467: begin  
rid<=0;
end
19'd171601: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=26;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6919;
 end   
19'd171602: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=96;
   mapp<=24;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10957;
 end   
19'd171603: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=39;
   mapp<=73;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12964;
 end   
19'd171604: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=85;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=10397;
 end   
19'd171605: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=74;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6428;
 end   
19'd171606: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=27;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6491;
 end   
19'd171607: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd171608: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd171609: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=68;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=13961;
 end   
19'd171610: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=18;
   mapp<=82;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=16957;
 end   
19'd171611: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=22;
   mapp<=15;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=16200;
 end   
19'd171612: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=7;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=13023;
 end   
19'd171613: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=95;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=14700;
 end   
19'd171614: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=20;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=10711;
 end   
19'd171615: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd171616: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd171617: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd171759: begin  
rid<=1;
end
19'd171760: begin  
end
19'd171761: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd171762: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd171763: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd171764: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd171765: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd171766: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd171767: begin  
rid<=0;
end
19'd171901: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=66;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8873;
 end   
19'd171902: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=89;
   mapp<=73;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9784;
 end   
19'd171903: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=90;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9611;
 end   
19'd171904: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=87;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5571;
 end   
19'd171905: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=33;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=8017;
 end   
19'd171906: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=93;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7924;
 end   
19'd171907: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=62;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=2876;
 end   
19'd171908: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=8;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=3789;
 end   
19'd171909: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=47;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd171910: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=92;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=9429;
 end   
19'd171911: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=2;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=14258;
 end   
19'd171912: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=93;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=12764;
 end   
19'd171913: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=56;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=8731;
 end   
19'd171914: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=60;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=12973;
 end   
19'd171915: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=97;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=10425;
 end   
19'd171916: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=42;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=5006;
 end   
19'd171917: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=40;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=4949;
 end   
19'd171918: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=20;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd171919: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd172061: begin  
rid<=1;
end
19'd172062: begin  
end
19'd172063: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd172064: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd172065: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd172066: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd172067: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd172068: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd172069: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd172070: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd172071: begin  
rid<=0;
end
19'd172201: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=17;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=15108;
 end   
19'd172202: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=53;
   mapp<=17;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=21029;
 end   
19'd172203: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=26;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd172204: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=7;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd172205: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=30;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd172206: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=68;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd172207: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=44;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd172208: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=87;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd172209: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=8;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd172210: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd172211: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=40;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=32702;
 end   
19'd172212: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=50;
   mapp<=30;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=38312;
 end   
19'd172213: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=15;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd172214: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=61;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd172215: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=51;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd172216: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=55;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd172217: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=3;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd172218: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=68;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd172219: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=41;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd172220: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd172221: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd172363: begin  
rid<=1;
end
19'd172364: begin  
end
19'd172365: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd172366: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd172367: begin  
rid<=0;
end
19'd172501: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=58;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=30460;
 end   
19'd172502: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=28;
   mapp<=78;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=28964;
 end   
19'd172503: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=45;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd172504: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=56;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd172505: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=84;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd172506: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=41;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd172507: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=32;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd172508: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=16;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd172509: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=59;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd172510: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=67;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd172511: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd172512: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=27;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=58090;
 end   
19'd172513: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=17;
   mapp<=66;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=54738;
 end   
19'd172514: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=85;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd172515: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=98;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd172516: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=25;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd172517: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=65;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd172518: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=96;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd172519: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=47;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd172520: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd172521: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=97;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd172522: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd172523: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd172665: begin  
rid<=1;
end
19'd172666: begin  
end
19'd172667: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd172668: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd172669: begin  
rid<=0;
end
19'd172801: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=51;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12192;
 end   
19'd172802: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=22;
   mapp<=57;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10658;
 end   
19'd172803: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=71;
   mapp<=68;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7978;
 end   
19'd172804: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=86;
   mapp<=27;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=8096;
 end   
19'd172805: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=58;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd172806: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=74;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd172807: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd172808: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd172809: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd172810: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=14;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=38468;
 end   
19'd172811: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=64;
   mapp<=94;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=29981;
 end   
19'd172812: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=65;
   mapp<=66;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=25207;
 end   
19'd172813: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=28;
   mapp<=21;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=33877;
 end   
19'd172814: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=98;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd172815: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=71;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd172816: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd172817: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd172818: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd172819: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd172961: begin  
rid<=1;
end
19'd172962: begin  
end
19'd172963: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd172964: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd172965: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd172966: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd172967: begin  
rid<=0;
end
19'd173101: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9407;
 end   
19'd173102: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=69;
   mapp<=41;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11344;
 end   
19'd173103: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=10;
   mapp<=19;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8214;
 end   
19'd173104: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=47;
   mapp<=47;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=14217;
 end   
19'd173105: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=14;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd173106: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=77;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd173107: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=63;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd173108: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=22;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd173109: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=95;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd173110: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=52;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd173111: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=74;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=26247;
 end   
19'd173112: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=18;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18350;
 end   
19'd173113: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=83;
   mapp<=83;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=16969;
 end   
19'd173114: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=3;
   mapp<=17;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=21136;
 end   
19'd173115: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=31;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd173116: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=61;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd173117: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=65;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd173118: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=3;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd173119: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=1;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd173120: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=45;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd173121: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd173263: begin  
rid<=1;
end
19'd173264: begin  
end
19'd173265: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd173266: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd173267: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd173268: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd173269: begin  
rid<=0;
end
19'd173401: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=95;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=31614;
 end   
19'd173402: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=88;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=26395;
 end   
19'd173403: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=31;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd173404: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=48;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd173405: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=85;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd173406: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=48;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd173407: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=54;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd173408: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=95;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd173409: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=34;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd173410: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=52;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd173411: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=68;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd173412: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=43;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=50440;
 end   
19'd173413: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=30;
   mapp<=9;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=45300;
 end   
19'd173414: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=33;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd173415: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=89;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd173416: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=10;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd173417: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=37;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd173418: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=12;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd173419: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=45;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd173420: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=8;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd173421: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=46;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd173422: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=60;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd173423: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd173565: begin  
rid<=1;
end
19'd173566: begin  
end
19'd173567: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd173568: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd173569: begin  
rid<=0;
end
19'd173701: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=24;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5682;
 end   
19'd173702: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=20;
   mapp<=75;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8042;
 end   
19'd173703: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=86;
   mapp<=45;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10510;
 end   
19'd173704: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=62;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=10298;
 end   
19'd173705: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=95;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4350;
 end   
19'd173706: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=80;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=5166;
 end   
19'd173707: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=5;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=7694;
 end   
19'd173708: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd173709: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd173710: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=56;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14103;
 end   
19'd173711: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=79;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=14602;
 end   
19'd173712: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=5;
   mapp<=32;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=16821;
 end   
19'd173713: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=56;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=15295;
 end   
19'd173714: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=19;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=11267;
 end   
19'd173715: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=72;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=12275;
 end   
19'd173716: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=33;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=16983;
 end   
19'd173717: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd173718: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd173719: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd173861: begin  
rid<=1;
end
19'd173862: begin  
end
19'd173863: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd173864: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd173865: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd173866: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd173867: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd173868: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd173869: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd173870: begin  
rid<=0;
end
19'd174001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=23;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=782;
 end   
19'd174002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=60;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1390;
 end   
19'd174003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=69;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1607;
 end   
19'd174004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=28;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=674;
 end   
19'd174005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=93;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2179;
 end   
19'd174006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=63;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=1499;
 end   
19'd174007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=35;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=865;
 end   
19'd174008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=22;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=576;
 end   
19'd174009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=91;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=2173;
 end   
19'd174010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=13;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=389;
 end   
19'd174011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=73;
   pp<=100;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[10]<=1779;
 end   
19'd174012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=58;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=1188;
 end   
19'd174013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=66;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=5218;
 end   
19'd174014: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=80;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=6247;
 end   
19'd174015: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=62;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=4270;
 end   
19'd174016: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=66;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=6007;
 end   
19'd174017: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=27;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=3065;
 end   
19'd174018: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=59;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=4287;
 end   
19'd174019: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=19;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=1678;
 end   
19'd174020: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=9;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=2695;
 end   
19'd174021: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=76;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=4797;
 end   
19'd174022: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=28;
   pp<=100;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[10]<=3403;
 end   
19'd174023: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd174165: begin  
rid<=1;
end
19'd174166: begin  
end
19'd174167: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd174168: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd174169: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd174170: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd174171: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd174172: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd174173: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd174174: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd174175: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd174176: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd174177: begin  
check0<=expctdoutput[10]-outcheck0;
end
19'd174178: begin  
rid<=0;
end
19'd174301: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=92;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16857;
 end   
19'd174302: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=15;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=20135;
 end   
19'd174303: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=99;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd174304: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=67;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd174305: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=58;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd174306: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd174307: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=83;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=26139;
 end   
19'd174308: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=89;
   mapp<=20;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=30877;
 end   
19'd174309: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=34;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd174310: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=27;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd174311: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=25;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd174312: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd174313: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd174455: begin  
rid<=1;
end
19'd174456: begin  
end
19'd174457: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd174458: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd174459: begin  
rid<=0;
end
19'd174601: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=52;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2049;
 end   
19'd174602: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=19;
   mapp<=23;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1282;
 end   
19'd174603: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=4;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2071;
 end   
19'd174604: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=97;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6062;
 end   
19'd174605: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=52;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4511;
 end   
19'd174606: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=93;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=5950;
 end   
19'd174607: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=56;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=3428;
 end   
19'd174608: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=24;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=2648;
 end   
19'd174609: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=70;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=4518;
 end   
19'd174610: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd174611: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=81;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=11706;
 end   
19'd174612: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=33;
   mapp<=57;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8209;
 end   
19'd174613: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=10018;
 end   
19'd174614: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=69;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=14918;
 end   
19'd174615: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=99;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=15071;
 end   
19'd174616: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=77;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=13111;
 end   
19'd174617: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=28;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=7214;
 end   
19'd174618: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=46;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=7892;
 end   
19'd174619: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=46;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=10653;
 end   
19'd174620: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd174621: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd174763: begin  
rid<=1;
end
19'd174764: begin  
end
19'd174765: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd174766: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd174767: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd174768: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd174769: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd174770: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd174771: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd174772: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd174773: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd174774: begin  
rid<=0;
end
19'd174901: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=38;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=19905;
 end   
19'd174902: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=39;
   mapp<=44;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=18622;
 end   
19'd174903: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=92;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd174904: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=14;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd174905: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=29;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd174906: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=60;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd174907: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=68;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd174908: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=52;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=37130;
 end   
19'd174909: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=69;
   mapp<=37;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=35172;
 end   
19'd174910: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=22;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd174911: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=71;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd174912: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=48;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd174913: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=96;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd174914: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=36;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd174915: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd175057: begin  
rid<=1;
end
19'd175058: begin  
end
19'd175059: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd175060: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd175061: begin  
rid<=0;
end
19'd175201: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=86;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16888;
 end   
19'd175202: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=45;
   mapp<=8;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=20593;
 end   
19'd175203: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=70;
   mapp<=91;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=25564;
 end   
19'd175204: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=13;
   mapp<=21;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=20820;
 end   
19'd175205: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=48;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd175206: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=79;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd175207: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=86;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd175208: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=1;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd175209: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd175210: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd175211: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd175212: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=84;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=40426;
 end   
19'd175213: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=35;
   mapp<=14;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=41224;
 end   
19'd175214: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=89;
   mapp<=65;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=47570;
 end   
19'd175215: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=91;
   mapp<=23;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=42439;
 end   
19'd175216: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=36;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd175217: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=2;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd175218: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=74;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd175219: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=86;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd175220: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd175221: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd175222: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd175223: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd175365: begin  
rid<=1;
end
19'd175366: begin  
end
19'd175367: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd175368: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd175369: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd175370: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd175371: begin  
rid<=0;
end
19'd175501: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=35;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=19289;
 end   
19'd175502: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=90;
   mapp<=31;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=27952;
 end   
19'd175503: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=78;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd175504: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=68;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd175505: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=19;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd175506: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd175507: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=65;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd175508: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=43;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd175509: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=69;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd175510: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=82;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd175511: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=80;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=41480;
 end   
19'd175512: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=6;
   mapp<=55;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=49645;
 end   
19'd175513: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=76;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd175514: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=86;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd175515: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=84;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd175516: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=23;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd175517: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=28;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd175518: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=27;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd175519: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=35;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd175520: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=32;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd175521: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd175663: begin  
rid<=1;
end
19'd175664: begin  
end
19'd175665: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd175666: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd175667: begin  
rid<=0;
end
19'd175801: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=36;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12134;
 end   
19'd175802: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=66;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12913;
 end   
19'd175803: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=10;
   mapp<=31;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=16570;
 end   
19'd175804: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=22;
   mapp<=62;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=10605;
 end   
19'd175805: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=59;
   mapp<=2;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=11422;
 end   
19'd175806: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=26;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd175807: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=44;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd175808: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd175809: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd175810: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd175811: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd175812: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=5;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=25369;
 end   
19'd175813: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=97;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=29738;
 end   
19'd175814: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=31;
   mapp<=46;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=38782;
 end   
19'd175815: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=78;
   mapp<=44;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=26069;
 end   
19'd175816: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=23;
   mapp<=36;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=35772;
 end   
19'd175817: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=61;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd175818: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=60;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd175819: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd175820: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd175821: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd175822: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd175823: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd175965: begin  
rid<=1;
end
19'd175966: begin  
end
19'd175967: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd175968: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd175969: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd175970: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd175971: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd175972: begin  
rid<=0;
end
19'd176101: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=51;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=18419;
 end   
19'd176102: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=83;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd176103: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=78;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd176104: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=18;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd176105: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=25;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd176106: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=42;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd176107: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=62;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=35757;
 end   
19'd176108: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=55;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd176109: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=91;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd176110: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=70;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd176111: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=7;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd176112: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=90;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd176113: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd176255: begin  
rid<=1;
end
19'd176256: begin  
end
19'd176257: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd176258: begin  
rid<=0;
end
19'd176401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=30;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=17438;
 end   
19'd176402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=1;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd176403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=86;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd176404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=33;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd176405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=73;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd176406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=46;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd176407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=15;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd176408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=81;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd176409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=87;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=50781;
 end   
19'd176410: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=80;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd176411: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=55;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd176412: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=43;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd176413: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=99;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd176414: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=43;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd176415: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=15;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd176416: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=79;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd176417: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd176559: begin  
rid<=1;
end
19'd176560: begin  
end
19'd176561: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd176562: begin  
rid<=0;
end
19'd176701: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=17;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1156;
 end   
19'd176702: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=18;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1234;
 end   
19'd176703: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=76;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5188;
 end   
19'd176704: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=19;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1322;
 end   
19'd176705: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=81;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5548;
 end   
19'd176706: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=18;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=1274;
 end   
19'd176707: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=17;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=1216;
 end   
19'd176708: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=80;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7396;
 end   
19'd176709: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=57;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=5680;
 end   
19'd176710: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=76;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=11116;
 end   
19'd176711: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=43;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=4676;
 end   
19'd176712: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=29;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=7810;
 end   
19'd176713: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=36;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=4082;
 end   
19'd176714: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=10;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=1996;
 end   
19'd176715: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd176857: begin  
rid<=1;
end
19'd176858: begin  
end
19'd176859: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd176860: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd176861: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd176862: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd176863: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd176864: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd176865: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd176866: begin  
rid<=0;
end
19'd177001: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=4;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10663;
 end   
19'd177002: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=58;
   mapp<=7;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12930;
 end   
19'd177003: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=83;
   mapp<=79;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8627;
 end   
19'd177004: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=38;
   mapp<=96;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5290;
 end   
19'd177005: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=9;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5265;
 end   
19'd177006: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=52;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7617;
 end   
19'd177007: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd177008: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd177009: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd177010: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=69;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=20725;
 end   
19'd177011: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=84;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=25143;
 end   
19'd177012: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=90;
   mapp<=11;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=20912;
 end   
19'd177013: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=6;
   mapp<=49;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=22831;
 end   
19'd177014: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=77;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=25080;
 end   
19'd177015: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=80;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=26529;
 end   
19'd177016: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd177017: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd177018: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd177019: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd177161: begin  
rid<=1;
end
19'd177162: begin  
end
19'd177163: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd177164: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd177165: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd177166: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd177167: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd177168: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd177169: begin  
rid<=0;
end
19'd177301: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=27;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=28012;
 end   
19'd177302: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=95;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=29916;
 end   
19'd177303: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=87;
   mapp<=48;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=28417;
 end   
19'd177304: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=63;
   mapp<=33;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=25076;
 end   
19'd177305: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=62;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd177306: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=93;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd177307: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=53;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd177308: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=14;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd177309: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=85;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd177310: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=57;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd177311: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=2;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd177312: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=90;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=56444;
 end   
19'd177313: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=20;
   mapp<=23;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=52121;
 end   
19'd177314: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=48;
   mapp<=39;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=47992;
 end   
19'd177315: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=39;
   mapp<=23;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=46877;
 end   
19'd177316: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=6;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd177317: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=60;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd177318: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=54;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd177319: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=99;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd177320: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=9;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd177321: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=3;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd177322: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=54;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd177323: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd177465: begin  
rid<=1;
end
19'd177466: begin  
end
19'd177467: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd177468: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd177469: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd177470: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd177471: begin  
rid<=0;
end
19'd177601: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=7;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4890;
 end   
19'd177602: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=30;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7071;
 end   
19'd177603: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=47;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd177604: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=48;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd177605: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=80;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17876;
 end   
19'd177606: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=37;
   mapp<=98;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18774;
 end   
19'd177607: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=32;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd177608: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=80;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd177609: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd177751: begin  
rid<=1;
end
19'd177752: begin  
end
19'd177753: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd177754: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd177755: begin  
rid<=0;
end
19'd177901: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=65;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1365;
 end   
19'd177902: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=84;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1774;
 end   
19'd177903: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=73;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1553;
 end   
19'd177904: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=59;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1269;
 end   
19'd177905: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=30;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=670;
 end   
19'd177906: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=34;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=764;
 end   
19'd177907: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=36;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=816;
 end   
19'd177908: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=10;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=2305;
 end   
19'd177909: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=19;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=3560;
 end   
19'd177910: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=10;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=2493;
 end   
19'd177911: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=69;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=7755;
 end   
19'd177912: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=89;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=9036;
 end   
19'd177913: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=34;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=3960;
 end   
19'd177914: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=85;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=8806;
 end   
19'd177915: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd178057: begin  
rid<=1;
end
19'd178058: begin  
end
19'd178059: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd178060: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd178061: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd178062: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd178063: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd178064: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd178065: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd178066: begin  
rid<=0;
end
19'd178201: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=16;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14729;
 end   
19'd178202: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=93;
   mapp<=54;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=14954;
 end   
19'd178203: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=38;
   mapp<=67;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12948;
 end   
19'd178204: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=95;
   mapp<=52;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=11617;
 end   
19'd178205: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=71;
   mapp<=11;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=21606;
 end   
19'd178206: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd178207: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd178208: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd178209: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd178210: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=10;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17587;
 end   
19'd178211: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=11;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=17877;
 end   
19'd178212: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=17;
   mapp<=35;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15531;
 end   
19'd178213: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=14;
   mapp<=27;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=14290;
 end   
19'd178214: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=17;
   mapp<=44;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=25236;
 end   
19'd178215: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd178216: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd178217: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd178218: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd178219: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd178361: begin  
rid<=1;
end
19'd178362: begin  
end
19'd178363: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd178364: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd178365: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd178366: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd178367: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd178368: begin  
rid<=0;
end
19'd178501: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=77;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=18144;
 end   
19'd178502: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=61;
   mapp<=90;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8780;
 end   
19'd178503: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=9;
   mapp<=4;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=18419;
 end   
19'd178504: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=96;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd178505: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=44;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd178506: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=19;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd178507: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd178508: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=56;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=26073;
 end   
19'd178509: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=74;
   mapp<=63;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20859;
 end   
19'd178510: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=4;
   mapp<=79;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=29721;
 end   
19'd178511: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=74;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd178512: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=3;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd178513: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd178514: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd178515: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd178657: begin  
rid<=1;
end
19'd178658: begin  
end
19'd178659: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd178660: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd178661: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd178662: begin  
rid<=0;
end
19'd178801: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=53;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10204;
 end   
19'd178802: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=47;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12862;
 end   
19'd178803: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=21;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd178804: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=39;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd178805: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=39;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd178806: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=19;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd178807: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=25;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd178808: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=59;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd178809: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=92;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd178810: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=49;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=30860;
 end   
19'd178811: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=45;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=32870;
 end   
19'd178812: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=62;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd178813: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=28;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd178814: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=88;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd178815: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=84;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd178816: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=31;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd178817: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=43;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd178818: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=60;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd178819: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd178961: begin  
rid<=1;
end
19'd178962: begin  
end
19'd178963: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd178964: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd178965: begin  
rid<=0;
end
19'd179101: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=32;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3504;
 end   
19'd179102: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=52;
   mapp<=12;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4798;
 end   
19'd179103: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=9;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=986;
 end   
19'd179104: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=13;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1512;
 end   
19'd179105: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=26;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2812;
 end   
19'd179106: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=36;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=3350;
 end   
19'd179107: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=5;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=630;
 end   
19'd179108: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=10;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=1918;
 end   
19'd179109: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=79;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=7574;
 end   
19'd179110: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=32;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd179111: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=3;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=4770;
 end   
19'd179112: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=30;
   mapp<=36;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8026;
 end   
19'd179113: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=38;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=3450;
 end   
19'd179114: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=3;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=4938;
 end   
19'd179115: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=90;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=11920;
 end   
19'd179116: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=98;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=12990;
 end   
19'd179117: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=99;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=9000;
 end   
19'd179118: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=62;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=7418;
 end   
19'd179119: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=46;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=13882;
 end   
19'd179120: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=96;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd179121: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd179263: begin  
rid<=1;
end
19'd179264: begin  
end
19'd179265: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd179266: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd179267: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd179268: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd179269: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd179270: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd179271: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd179272: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd179273: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd179274: begin  
rid<=0;
end
19'd179401: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=67;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=18955;
 end   
19'd179402: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=76;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=16034;
 end   
19'd179403: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=34;
   mapp<=38;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11848;
 end   
19'd179404: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=56;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd179405: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=65;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd179406: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=15;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd179407: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=22;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd179408: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=81;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=29172;
 end   
19'd179409: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=56;
   mapp<=86;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=26020;
 end   
19'd179410: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=49;
   mapp<=7;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=20442;
 end   
19'd179411: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=25;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd179412: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=53;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd179413: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=52;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd179414: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd179415: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd179557: begin  
rid<=1;
end
19'd179558: begin  
end
19'd179559: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd179560: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd179561: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd179562: begin  
rid<=0;
end
19'd179701: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=60;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2654;
 end   
19'd179702: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=11;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd179703: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=44;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7418;
 end   
19'd179704: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=20;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd179705: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd179847: begin  
rid<=1;
end
19'd179848: begin  
end
19'd179849: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd179850: begin  
rid<=0;
end
19'd180001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=49;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=26625;
 end   
19'd180002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=16;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd180003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=60;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd180004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=11;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd180005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=32;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd180006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=82;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd180007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=38;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd180008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=84;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd180009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=59;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd180010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=68;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd180011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=89;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd180012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=47;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=44575;
 end   
19'd180013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=33;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd180014: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=79;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd180015: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=32;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd180016: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=5;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd180017: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=32;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd180018: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=47;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd180019: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=13;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd180020: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=9;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd180021: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=30;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd180022: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=57;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd180023: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd180165: begin  
rid<=1;
end
19'd180166: begin  
end
19'd180167: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd180168: begin  
rid<=0;
end
19'd180301: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=40;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=21787;
 end   
19'd180302: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=88;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=21062;
 end   
19'd180303: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=55;
   mapp<=26;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=23962;
 end   
19'd180304: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=71;
   mapp<=81;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=25118;
 end   
19'd180305: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=70;
   mapp<=69;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=20358;
 end   
19'd180306: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=79;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=18841;
 end   
19'd180307: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd180308: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd180309: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd180310: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd180311: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=40;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=31153;
 end   
19'd180312: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=7;
   mapp<=79;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=29365;
 end   
19'd180313: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=91;
   mapp<=28;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=30624;
 end   
19'd180314: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=11;
   mapp<=3;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=34622;
 end   
19'd180315: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=98;
   mapp<=24;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=27163;
 end   
19'd180316: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=45;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=33309;
 end   
19'd180317: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd180318: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd180319: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd180320: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd180321: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd180463: begin  
rid<=1;
end
19'd180464: begin  
end
19'd180465: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd180466: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd180467: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd180468: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd180469: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd180470: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd180471: begin  
rid<=0;
end
19'd180601: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=7;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6030;
 end   
19'd180602: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=41;
   mapp<=15;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4694;
 end   
19'd180603: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=13;
   mapp<=10;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4294;
 end   
19'd180604: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=94;
   mapp<=26;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7084;
 end   
19'd180605: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=81;
   mapp<=33;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5590;
 end   
19'd180606: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=9;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6822;
 end   
19'd180607: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=23;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=7945;
 end   
19'd180608: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd180609: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd180610: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd180611: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd180612: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=41;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=15437;
 end   
19'd180613: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=44;
   mapp<=50;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12898;
 end   
19'd180614: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=19;
   mapp<=96;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=13406;
 end   
19'd180615: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=24;
   mapp<=71;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=15491;
 end   
19'd180616: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=49;
   mapp<=14;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=9611;
 end   
19'd180617: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=5;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=13657;
 end   
19'd180618: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=34;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=18629;
 end   
19'd180619: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd180620: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd180621: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd180622: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd180623: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd180765: begin  
rid<=1;
end
19'd180766: begin  
end
19'd180767: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd180768: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd180769: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd180770: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd180771: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd180772: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd180773: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd180774: begin  
rid<=0;
end
19'd180901: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=82;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8744;
 end   
19'd180902: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=78;
   mapp<=69;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3415;
 end   
19'd180903: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=3;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2903;
 end   
19'd180904: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=40;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3947;
 end   
19'd180905: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=33;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2911;
 end   
19'd180906: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=22;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6817;
 end   
19'd180907: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=85;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd180908: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=80;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=11704;
 end   
19'd180909: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=16;
   mapp<=75;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=6017;
 end   
19'd180910: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=30;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=4763;
 end   
19'd180911: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=16;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=8349;
 end   
19'd180912: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=54;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=7399;
 end   
19'd180913: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=44;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=14385;
 end   
19'd180914: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd180915: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd181057: begin  
rid<=1;
end
19'd181058: begin  
end
19'd181059: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd181060: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd181061: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd181062: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd181063: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd181064: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd181065: begin  
rid<=0;
end
19'd181201: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=57;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5163;
 end   
19'd181202: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=46;
   mapp<=54;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5844;
 end   
19'd181203: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=68;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4242;
 end   
19'd181204: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=19;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd181205: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=11631;
 end   
19'd181206: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=84;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12060;
 end   
19'd181207: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=36;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=6334;
 end   
19'd181208: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=8;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd181209: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd181351: begin  
rid<=1;
end
19'd181352: begin  
end
19'd181353: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd181354: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd181355: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd181356: begin  
rid<=0;
end
19'd181501: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=47;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16084;
 end   
19'd181502: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=65;
   mapp<=89;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=16704;
 end   
19'd181503: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=72;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd181504: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=4;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd181505: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=35;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd181506: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=83;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd181507: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=28;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd181508: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=30;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd181509: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd181510: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=19;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=40755;
 end   
19'd181511: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=28;
   mapp<=29;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=39113;
 end   
19'd181512: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=51;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd181513: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=75;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd181514: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=61;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd181515: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=97;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd181516: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=50;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd181517: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=19;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd181518: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd181519: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd181661: begin  
rid<=1;
end
19'd181662: begin  
end
19'd181663: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd181664: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd181665: begin  
rid<=0;
end
19'd181801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=15;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1935;
 end   
19'd181802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=24;
   mapp<=30;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3694;
 end   
19'd181803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=58;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd181804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=40;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7355;
 end   
19'd181805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=73;
   mapp<=20;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12561;
 end   
19'd181806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=82;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd181807: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd181949: begin  
rid<=1;
end
19'd181950: begin  
end
19'd181951: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd181952: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd181953: begin  
rid<=0;
end
19'd182101: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=61;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5761;
 end   
19'd182102: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=67;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5185;
 end   
19'd182103: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=80;
   mapp<=27;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7634;
 end   
19'd182104: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=46;
   mapp<=21;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=9227;
 end   
19'd182105: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=34;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=9356;
 end   
19'd182106: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=40;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6877;
 end   
19'd182107: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=53;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=8612;
 end   
19'd182108: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=7;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=9971;
 end   
19'd182109: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd182110: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd182111: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd182112: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=65;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=18398;
 end   
19'd182113: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=60;
   mapp<=85;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=19306;
 end   
19'd182114: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=26;
   mapp<=52;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15392;
 end   
19'd182115: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=70;
   mapp<=41;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=17666;
 end   
19'd182116: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=63;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=14813;
 end   
19'd182117: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=4;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=15563;
 end   
19'd182118: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=27;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=16207;
 end   
19'd182119: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=6;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=21029;
 end   
19'd182120: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd182121: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd182122: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd182123: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd182265: begin  
rid<=1;
end
19'd182266: begin  
end
19'd182267: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd182268: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd182269: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd182270: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd182271: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd182272: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd182273: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd182274: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd182275: begin  
rid<=0;
end
19'd182401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=95;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=21063;
 end   
19'd182402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=72;
   mapp<=57;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=19270;
 end   
19'd182403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=46;
   mapp<=69;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=21224;
 end   
19'd182404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=3;
   mapp<=31;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=18497;
 end   
19'd182405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=98;
   mapp<=99;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=21376;
 end   
19'd182406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=73;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=18277;
 end   
19'd182407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=78;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=18752;
 end   
19'd182408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd182409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd182410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd182411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd182412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=61;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=33690;
 end   
19'd182413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=40;
   mapp<=47;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=32053;
 end   
19'd182414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=68;
   mapp<=51;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=30693;
 end   
19'd182415: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=28;
   mapp<=84;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=30349;
 end   
19'd182416: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=46;
   mapp<=5;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=27909;
 end   
19'd182417: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=44;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=30457;
 end   
19'd182418: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=31;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=29577;
 end   
19'd182419: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd182420: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd182421: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd182422: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd182423: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd182565: begin  
rid<=1;
end
19'd182566: begin  
end
19'd182567: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd182568: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd182569: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd182570: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd182571: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd182572: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd182573: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd182574: begin  
rid<=0;
end
19'd182701: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=47;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12165;
 end   
19'd182702: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=66;
   mapp<=23;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=16375;
 end   
19'd182703: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=39;
   mapp<=75;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=13851;
 end   
19'd182704: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=86;
   mapp<=27;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=17122;
 end   
19'd182705: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=74;
   mapp<=12;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=16663;
 end   
19'd182706: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=57;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd182707: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=85;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd182708: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=47;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd182709: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=47;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd182710: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=20;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=20602;
 end   
19'd182711: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=56;
   mapp<=36;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=28972;
 end   
19'd182712: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=61;
   mapp<=68;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=21755;
 end   
19'd182713: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=93;
   mapp<=11;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=26913;
 end   
19'd182714: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=22;
   mapp<=25;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=20744;
 end   
19'd182715: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=75;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd182716: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=4;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd182717: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=24;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd182718: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=3;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd182719: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd182861: begin  
rid<=1;
end
19'd182862: begin  
end
19'd182863: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd182864: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd182865: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd182866: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd182867: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd182868: begin  
rid<=0;
end
19'd183001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=4;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9027;
 end   
19'd183002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=40;
   mapp<=30;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9151;
 end   
19'd183003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=73;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd183004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=22;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd183005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=31;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd183006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=82;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd183007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=55;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14663;
 end   
19'd183008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=24;
   mapp<=20;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=16493;
 end   
19'd183009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=34;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd183010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=18;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd183011: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=72;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd183012: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=56;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd183013: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd183155: begin  
rid<=1;
end
19'd183156: begin  
end
19'd183157: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd183158: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd183159: begin  
rid<=0;
end
19'd183301: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=15;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3690;
 end   
19'd183302: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=59;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5628;
 end   
19'd183303: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=56;
   mapp<=3;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6274;
 end   
19'd183304: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=72;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd183305: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=74;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd183306: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=15;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=10716;
 end   
19'd183307: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=59;
   mapp<=92;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=13675;
 end   
19'd183308: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=64;
   mapp<=17;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=10077;
 end   
19'd183309: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=9;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd183310: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=47;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd183311: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd183453: begin  
rid<=1;
end
19'd183454: begin  
end
19'd183455: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd183456: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd183457: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd183458: begin  
rid<=0;
end
19'd183601: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=91;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1270;
 end   
19'd183602: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=29;
   mapp<=3;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=519;
 end   
19'd183603: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=44;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=640;
 end   
19'd183604: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=16;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=493;
 end   
19'd183605: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=85;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1226;
 end   
19'd183606: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=27;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd183607: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=94;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5893;
 end   
19'd183608: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=39;
   mapp<=39;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=1962;
 end   
19'd183609: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=4;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=4165;
 end   
19'd183610: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=87;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=5977;
 end   
19'd183611: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=67;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=4022;
 end   
19'd183612: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=15;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd183613: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd183755: begin  
rid<=1;
end
19'd183756: begin  
end
19'd183757: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd183758: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd183759: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd183760: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd183761: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd183762: begin  
rid<=0;
end
19'd183901: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=91;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=22825;
 end   
19'd183902: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=25;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=13168;
 end   
19'd183903: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=91;
   mapp<=87;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=21906;
 end   
19'd183904: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=6;
   mapp<=14;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=10952;
 end   
19'd183905: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=42;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd183906: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=23;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd183907: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=17;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd183908: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=37;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd183909: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=75;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd183910: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=14;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd183911: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=6;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd183912: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=83;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=51879;
 end   
19'd183913: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=63;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=41620;
 end   
19'd183914: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=82;
   mapp<=96;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=50166;
 end   
19'd183915: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=43;
   mapp<=27;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=36077;
 end   
19'd183916: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=70;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd183917: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=21;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd183918: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=71;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd183919: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=97;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd183920: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=68;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd183921: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=40;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd183922: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=57;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd183923: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd184065: begin  
rid<=1;
end
19'd184066: begin  
end
19'd184067: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd184068: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd184069: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd184070: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd184071: begin  
rid<=0;
end
19'd184201: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=48;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10707;
 end   
19'd184202: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=76;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd184203: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=31;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd184204: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=74;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd184205: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=78;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd184206: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=67;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd184207: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=60;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd184208: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=49;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=28367;
 end   
19'd184209: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=22;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd184210: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=28;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd184211: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=60;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd184212: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=16;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd184213: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=67;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd184214: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=43;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd184215: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd184357: begin  
rid<=1;
end
19'd184358: begin  
end
19'd184359: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd184360: begin  
rid<=0;
end
19'd184501: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=19;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=23349;
 end   
19'd184502: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=43;
   mapp<=66;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=29541;
 end   
19'd184503: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=93;
   mapp<=23;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=21918;
 end   
19'd184504: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=46;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd184505: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=23;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd184506: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=77;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd184507: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=98;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd184508: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=32;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd184509: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=75;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd184510: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd184511: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd184512: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=28;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=41694;
 end   
19'd184513: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=41;
   mapp<=82;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=46514;
 end   
19'd184514: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=9;
   mapp<=96;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=38573;
 end   
19'd184515: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd184516: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=98;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd184517: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=17;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd184518: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=45;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd184519: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=27;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd184520: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=96;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd184521: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd184522: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd184523: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd184665: begin  
rid<=1;
end
19'd184666: begin  
end
19'd184667: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd184668: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd184669: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd184670: begin  
rid<=0;
end
19'd184801: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=71;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16328;
 end   
19'd184802: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=27;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10152;
 end   
19'd184803: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=92;
   mapp<=94;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11172;
 end   
19'd184804: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=49;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd184805: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=8;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd184806: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=85;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=28906;
 end   
19'd184807: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=52;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18112;
 end   
19'd184808: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=31;
   mapp<=19;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=17018;
 end   
19'd184809: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=36;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd184810: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=13;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd184811: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd184953: begin  
rid<=1;
end
19'd184954: begin  
end
19'd184955: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd184956: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd184957: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd184958: begin  
rid<=0;
end
19'd185101: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=50;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16982;
 end   
19'd185102: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=28;
   mapp<=13;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15963;
 end   
19'd185103: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=20;
   mapp<=55;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=14436;
 end   
19'd185104: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=32;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd185105: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=44;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd185106: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=18;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd185107: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=13;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd185108: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=91;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd185109: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd185110: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd185111: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=74;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=38357;
 end   
19'd185112: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=79;
   mapp<=51;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=42047;
 end   
19'd185113: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=28;
   mapp<=17;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=38417;
 end   
19'd185114: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=63;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd185115: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=79;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd185116: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=3;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd185117: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=52;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd185118: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=45;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd185119: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd185120: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd185121: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd185263: begin  
rid<=1;
end
19'd185264: begin  
end
19'd185265: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd185266: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd185267: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd185268: begin  
rid<=0;
end
19'd185401: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=99;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=15752;
 end   
19'd185402: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=92;
   mapp<=91;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11947;
 end   
19'd185403: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=50;
   mapp<=9;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7775;
 end   
19'd185404: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=42;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=14508;
 end   
19'd185405: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=60;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=18812;
 end   
19'd185406: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd185407: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd185408: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=10;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=24431;
 end   
19'd185409: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=54;
   mapp<=53;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=23304;
 end   
19'd185410: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=81;
   mapp<=67;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=18516;
 end   
19'd185411: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=89;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=20933;
 end   
19'd185412: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=65;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=23647;
 end   
19'd185413: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd185414: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd185415: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd185557: begin  
rid<=1;
end
19'd185558: begin  
end
19'd185559: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd185560: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd185561: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd185562: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd185563: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd185564: begin  
rid<=0;
end
19'd185701: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=66;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2772;
 end   
19'd185702: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=77;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3244;
 end   
19'd185703: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=47;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1994;
 end   
19'd185704: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=82;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3474;
 end   
19'd185705: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=7;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=334;
 end   
19'd185706: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=83;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=3536;
 end   
19'd185707: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=97;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=4134;
 end   
19'd185708: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=10;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=3732;
 end   
19'd185709: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=59;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8908;
 end   
19'd185710: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=80;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=9674;
 end   
19'd185711: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=7;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=4146;
 end   
19'd185712: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=33;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=3502;
 end   
19'd185713: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=59;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=9200;
 end   
19'd185714: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=86;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=12390;
 end   
19'd185715: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd185857: begin  
rid<=1;
end
19'd185858: begin  
end
19'd185859: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd185860: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd185861: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd185862: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd185863: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd185864: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd185865: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd185866: begin  
rid<=0;
end
19'd186001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=32;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=25137;
 end   
19'd186002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=46;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=23599;
 end   
19'd186003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=17;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd186004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=89;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd186005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=22;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd186006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=3;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd186007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=40;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd186008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=68;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd186009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=81;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd186010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=48;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd186011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd186012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=14;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=46649;
 end   
19'd186013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=23;
   mapp<=86;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=42807;
 end   
19'd186014: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=30;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd186015: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=95;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd186016: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=66;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd186017: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=41;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd186018: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=78;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd186019: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=42;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd186020: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=29;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd186021: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=14;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd186022: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd186023: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd186165: begin  
rid<=1;
end
19'd186166: begin  
end
19'd186167: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd186168: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd186169: begin  
rid<=0;
end
19'd186301: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=99;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8745;
 end   
19'd186302: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=15;
   mapp<=84;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4921;
 end   
19'd186303: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=43;
   mapp<=6;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6381;
 end   
19'd186304: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=34;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7792;
 end   
19'd186305: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=61;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6857;
 end   
19'd186306: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=26;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=4564;
 end   
19'd186307: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=30;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd186308: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd186309: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=98;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=27961;
 end   
19'd186310: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=94;
   mapp<=89;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=19312;
 end   
19'd186311: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=99;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=17905;
 end   
19'd186312: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=26;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=15787;
 end   
19'd186313: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=75;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=13083;
 end   
19'd186314: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=4;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=15093;
 end   
19'd186315: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=41;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd186316: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=96;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd186317: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd186459: begin  
rid<=1;
end
19'd186460: begin  
end
19'd186461: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd186462: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd186463: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd186464: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd186465: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd186466: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd186467: begin  
rid<=0;
end
19'd186601: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=7;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2593;
 end   
19'd186602: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=31;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd186603: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=43;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=6101;
 end   
19'd186604: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=24;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd186605: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd186747: begin  
rid<=1;
end
19'd186748: begin  
end
19'd186749: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd186750: begin  
rid<=0;
end
19'd186901: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=31;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10664;
 end   
19'd186902: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=90;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12508;
 end   
19'd186903: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=34;
   mapp<=23;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7874;
 end   
19'd186904: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=62;
   mapp<=12;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=11154;
 end   
19'd186905: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=18;
   mapp<=71;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=12723;
 end   
19'd186906: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=78;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=9115;
 end   
19'd186907: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=10;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=14706;
 end   
19'd186908: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=84;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd186909: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=69;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd186910: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=45;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd186911: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=81;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd186912: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=21;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14906;
 end   
19'd186913: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=60;
   mapp<=16;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=23574;
 end   
19'd186914: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=83;
   mapp<=4;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=17623;
 end   
19'd186915: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=13;
   mapp<=74;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=17288;
 end   
19'd186916: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=56;
   mapp<=1;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=20891;
 end   
19'd186917: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=22;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=18402;
 end   
19'd186918: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=53;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=25692;
 end   
19'd186919: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=32;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd186920: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=84;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd186921: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=71;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd186922: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=8;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd186923: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd187065: begin  
rid<=1;
end
19'd187066: begin  
end
19'd187067: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd187068: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd187069: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd187070: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd187071: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd187072: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd187073: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd187074: begin  
rid<=0;
end
19'd187201: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=58;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4350;
 end   
19'd187202: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=99;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7435;
 end   
19'd187203: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=59;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4445;
 end   
19'd187204: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=60;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4530;
 end   
19'd187205: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=37;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2815;
 end   
19'd187206: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=81;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6125;
 end   
19'd187207: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=55;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=4680;
 end   
19'd187208: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=38;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=7663;
 end   
19'd187209: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=39;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=4679;
 end   
19'd187210: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=12;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=4602;
 end   
19'd187211: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=55;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=3145;
 end   
19'd187212: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=97;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=6707;
 end   
19'd187213: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd187355: begin  
rid<=1;
end
19'd187356: begin  
end
19'd187357: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd187358: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd187359: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd187360: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd187361: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd187362: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd187363: begin  
rid<=0;
end
19'd187501: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=48;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14367;
 end   
19'd187502: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=5;
   mapp<=82;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=24610;
 end   
19'd187503: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=56;
   mapp<=28;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=24559;
 end   
19'd187504: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=53;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=29482;
 end   
19'd187505: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=65;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd187506: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=93;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd187507: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=85;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd187508: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=62;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd187509: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd187510: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd187511: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd187512: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=79;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=32248;
 end   
19'd187513: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=38;
   mapp<=16;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=46778;
 end   
19'd187514: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=46;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=51409;
 end   
19'd187515: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=72;
   mapp<=72;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=51818;
 end   
19'd187516: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=42;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd187517: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=4;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd187518: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=62;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd187519: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=36;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd187520: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd187521: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd187522: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd187523: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd187665: begin  
rid<=1;
end
19'd187666: begin  
end
19'd187667: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd187668: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd187669: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd187670: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd187671: begin  
rid<=0;
end
19'd187801: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=23;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2651;
 end   
19'd187802: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=73;
   mapp<=13;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3448;
 end   
19'd187803: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=43;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2177;
 end   
19'd187804: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=16;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3318;
 end   
19'd187805: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=40;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6946;
 end   
19'd187806: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=82;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=5002;
 end   
19'd187807: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=42;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=5844;
 end   
19'd187808: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=66;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=8523;
 end   
19'd187809: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd187810: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=61;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=9526;
 end   
19'd187811: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=93;
   mapp<=49;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12854;
 end   
19'd187812: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=69;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=13733;
 end   
19'd187813: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=79;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=12694;
 end   
19'd187814: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=49;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=12539;
 end   
19'd187815: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=28;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=6710;
 end   
19'd187816: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=13842;
 end   
19'd187817: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=86;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=21767;
 end   
19'd187818: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd187819: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd187961: begin  
rid<=1;
end
19'd187962: begin  
end
19'd187963: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd187964: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd187965: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd187966: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd187967: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd187968: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd187969: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd187970: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd187971: begin  
rid<=0;
end
19'd188101: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=39;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16720;
 end   
19'd188102: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=89;
   mapp<=47;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15186;
 end   
19'd188103: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=52;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=15441;
 end   
19'd188104: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=54;
   mapp<=44;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=18879;
 end   
19'd188105: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=96;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd188106: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=51;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd188107: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd188108: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd188109: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd188110: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=96;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=30402;
 end   
19'd188111: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=35;
   mapp<=75;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=31710;
 end   
19'd188112: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=61;
   mapp<=21;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=29504;
 end   
19'd188113: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=14;
   mapp<=67;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=35122;
 end   
19'd188114: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=54;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd188115: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=70;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd188116: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd188117: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd188118: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd188119: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd188261: begin  
rid<=1;
end
19'd188262: begin  
end
19'd188263: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd188264: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd188265: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd188266: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd188267: begin  
rid<=0;
end
19'd188401: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=96;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=15991;
 end   
19'd188402: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=23;
   mapp<=71;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12310;
 end   
19'd188403: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=56;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11490;
 end   
19'd188404: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=16;
   mapp<=30;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=9277;
 end   
19'd188405: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=90;
   mapp<=71;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=10936;
 end   
19'd188406: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd188407: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd188408: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd188409: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd188410: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=28;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=21904;
 end   
19'd188411: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=64;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=16380;
 end   
19'd188412: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=21;
   mapp<=23;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=14144;
 end   
19'd188413: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=9;
   mapp<=22;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=11492;
 end   
19'd188414: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=1;
   mapp<=8;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=14869;
 end   
19'd188415: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd188416: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd188417: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd188418: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd188419: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd188561: begin  
rid<=1;
end
19'd188562: begin  
end
19'd188563: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd188564: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd188565: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd188566: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd188567: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd188568: begin  
rid<=0;
end
19'd188701: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=98;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1470;
 end   
19'd188702: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=25;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=385;
 end   
19'd188703: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=34;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=530;
 end   
19'd188704: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=52;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=810;
 end   
19'd188705: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=0;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=1470;
 end   
19'd188706: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=8;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=665;
 end   
19'd188707: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=65;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=2805;
 end   
19'd188708: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=47;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=2455;
 end   
19'd188709: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd188851: begin  
rid<=1;
end
19'd188852: begin  
end
19'd188853: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd188854: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd188855: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd188856: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd188857: begin  
rid<=0;
end
19'd189001: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=57;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14953;
 end   
19'd189002: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=91;
   mapp<=60;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11485;
 end   
19'd189003: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=97;
   mapp<=82;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12523;
 end   
19'd189004: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=39;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=8653;
 end   
19'd189005: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=92;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=11486;
 end   
19'd189006: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=25;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd189007: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=91;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd189008: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=18325;
 end   
19'd189009: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=22;
   mapp<=96;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20129;
 end   
19'd189010: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=70;
   mapp<=18;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=23681;
 end   
19'd189011: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=91;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=18908;
 end   
19'd189012: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=84;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=19016;
 end   
19'd189013: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=56;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd189014: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=59;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd189015: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd189157: begin  
rid<=1;
end
19'd189158: begin  
end
19'd189159: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd189160: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd189161: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd189162: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd189163: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd189164: begin  
rid<=0;
end
19'd189301: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=9;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1233;
 end   
19'd189302: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=23;
   mapp<=45;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1887;
 end   
19'd189303: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=64;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=803;
 end   
19'd189304: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=9;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1744;
 end   
19'd189305: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=71;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2220;
 end   
19'd189306: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=67;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=1941;
 end   
19'd189307: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=56;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=2703;
 end   
19'd189308: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=93;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=2747;
 end   
19'd189309: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=80;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=2847;
 end   
19'd189310: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=89;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=1190;
 end   
19'd189311: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd189312: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=35;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=1913;
 end   
19'd189313: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=15;
   mapp<=43;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=4442;
 end   
19'd189314: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=4108;
 end   
19'd189315: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=57;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=4564;
 end   
19'd189316: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=55;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=4700;
 end   
19'd189317: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=37;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=4601;
 end   
19'd189318: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=91;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=7118;
 end   
19'd189319: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=82;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=6967;
 end   
19'd189320: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=90;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=7002;
 end   
19'd189321: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=67;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=4840;
 end   
19'd189322: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd189323: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd189465: begin  
rid<=1;
end
19'd189466: begin  
end
19'd189467: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd189468: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd189469: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd189470: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd189471: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd189472: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd189473: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd189474: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd189475: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd189476: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd189477: begin  
rid<=0;
end
19'd189601: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=3;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=33282;
 end   
19'd189602: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=45;
   mapp<=74;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=28448;
 end   
19'd189603: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=57;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd189604: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=16;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd189605: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=57;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd189606: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=37;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd189607: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=65;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd189608: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=73;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd189609: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=97;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd189610: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=48;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd189611: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd189612: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=29;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=45280;
 end   
19'd189613: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=9;
   mapp<=60;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=40866;
 end   
19'd189614: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=40;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd189615: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=64;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd189616: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=49;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd189617: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=46;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd189618: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd189619: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=29;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd189620: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=58;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd189621: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=2;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd189622: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd189623: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd189765: begin  
rid<=1;
end
19'd189766: begin  
end
19'd189767: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd189768: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd189769: begin  
rid<=0;
end
19'd189901: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=66;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5325;
 end   
19'd189902: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=53;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9964;
 end   
19'd189903: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=72;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6309;
 end   
19'd189904: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=29;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3746;
 end   
19'd189905: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd189906: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=1;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=10172;
 end   
19'd189907: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=94;
   mapp<=51;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=13681;
 end   
19'd189908: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=39;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=13398;
 end   
19'd189909: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=75;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=11999;
 end   
19'd189910: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd189911: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd190053: begin  
rid<=1;
end
19'd190054: begin  
end
19'd190055: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd190056: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd190057: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd190058: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd190059: begin  
rid<=0;
end
19'd190201: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=1;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5682;
 end   
19'd190202: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=55;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7597;
 end   
19'd190203: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=61;
   mapp<=28;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5945;
 end   
19'd190204: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=23;
   mapp<=26;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5912;
 end   
19'd190205: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=78;
   mapp<=9;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5382;
 end   
19'd190206: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=13;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd190207: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=25;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd190208: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd190209: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=42;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd190210: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=34;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17004;
 end   
19'd190211: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=15;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=21900;
 end   
19'd190212: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=95;
   mapp<=65;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=18687;
 end   
19'd190213: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=35;
   mapp<=4;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=17178;
 end   
19'd190214: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=42;
   mapp<=41;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=17959;
 end   
19'd190215: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=75;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd190216: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=27;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd190217: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=17;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd190218: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=49;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd190219: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd190361: begin  
rid<=1;
end
19'd190362: begin  
end
19'd190363: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd190364: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd190365: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd190366: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd190367: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd190368: begin  
rid<=0;
end
19'd190501: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=49;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11101;
 end   
19'd190502: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=62;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=16287;
 end   
19'd190503: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=64;
   mapp<=27;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=13988;
 end   
19'd190504: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=43;
   mapp<=24;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7365;
 end   
19'd190505: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=11;
   mapp<=71;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=13336;
 end   
19'd190506: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=12;
   mapp<=82;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=17328;
 end   
19'd190507: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=86;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd190508: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=28;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd190509: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd190510: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=96;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd190511: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd190512: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=53;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=24934;
 end   
19'd190513: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=48;
   mapp<=31;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=30548;
 end   
19'd190514: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=99;
   mapp<=27;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=30221;
 end   
19'd190515: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=12;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=16000;
 end   
19'd190516: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=41;
   mapp<=30;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=27386;
 end   
19'd190517: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=54;
   mapp<=68;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=30167;
 end   
19'd190518: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd190519: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=51;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd190520: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=52;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd190521: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=68;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd190522: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=26;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd190523: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd190665: begin  
rid<=1;
end
19'd190666: begin  
end
19'd190667: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd190668: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd190669: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd190670: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd190671: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd190672: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd190673: begin  
rid<=0;
end
19'd190801: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=28;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=23485;
 end   
19'd190802: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=89;
   mapp<=21;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=28586;
 end   
19'd190803: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=28;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd190804: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=83;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd190805: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=85;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd190806: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=36;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd190807: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=23;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd190808: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=65;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd190809: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=76;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd190810: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd190811: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd190812: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=33;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=62011;
 end   
19'd190813: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=41;
   mapp<=78;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=68045;
 end   
19'd190814: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=76;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd190815: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=72;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd190816: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=48;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd190817: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=75;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd190818: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=12;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd190819: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=97;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd190820: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=93;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd190821: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=96;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd190822: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd190823: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd190965: begin  
rid<=1;
end
19'd190966: begin  
end
19'd190967: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd190968: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd190969: begin  
rid<=0;
end
19'd191101: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=45;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2790;
 end   
19'd191102: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=67;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4164;
 end   
19'd191103: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=26;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1632;
 end   
19'd191104: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=0;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=2790;
 end   
19'd191105: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=65;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=5789;
 end   
19'd191106: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=79;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=3607;
 end   
19'd191107: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd191249: begin  
rid<=1;
end
19'd191250: begin  
end
19'd191251: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd191252: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd191253: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd191254: begin  
rid<=0;
end
19'd191401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=21;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=17520;
 end   
19'd191402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=16;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=16456;
 end   
19'd191403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=15;
   mapp<=26;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=18100;
 end   
19'd191404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=60;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd191405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=29;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd191406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=66;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd191407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=83;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd191408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=8;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd191409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=5;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd191410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd191411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd191412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=19;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=37095;
 end   
19'd191413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=32;
   mapp<=69;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=39515;
 end   
19'd191414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=92;
   mapp<=44;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=41296;
 end   
19'd191415: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=2;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd191416: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=17;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd191417: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=26;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd191418: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=60;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd191419: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=11;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd191420: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=87;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd191421: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd191422: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd191423: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd191565: begin  
rid<=1;
end
19'd191566: begin  
end
19'd191567: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd191568: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd191569: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd191570: begin  
rid<=0;
end
19'd191701: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=10;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4691;
 end   
19'd191702: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=75;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2409;
 end   
19'd191703: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=9;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd191704: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd191705: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=81;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12920;
 end   
19'd191706: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=30;
   mapp<=73;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12842;
 end   
19'd191707: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=40;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd191708: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd191709: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd191851: begin  
rid<=1;
end
19'd191852: begin  
end
19'd191853: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd191854: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd191855: begin  
rid<=0;
end
19'd192001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=47;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5917;
 end   
19'd192002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=66;
   mapp<=9;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2308;
 end   
19'd192003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=6;
   mapp<=14;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5801;
 end   
19'd192004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=25;
   mapp<=46;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5836;
 end   
19'd192005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=27;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=7927;
 end   
19'd192006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=77;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=9853;
 end   
19'd192007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=56;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=8538;
 end   
19'd192008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=48;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=9800;
 end   
19'd192009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd192010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd192011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd192012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=18;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14611;
 end   
19'd192013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=12;
   mapp<=54;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=13762;
 end   
19'd192014: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=88;
   mapp<=24;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=16605;
 end   
19'd192015: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=74;
   mapp<=78;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=18954;
 end   
19'd192016: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=45;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=21459;
 end   
19'd192017: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=74;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=26303;
 end   
19'd192018: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=63;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=19098;
 end   
19'd192019: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=85;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=17224;
 end   
19'd192020: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd192021: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd192022: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd192023: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd192165: begin  
rid<=1;
end
19'd192166: begin  
end
19'd192167: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd192168: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd192169: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd192170: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd192171: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd192172: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd192173: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd192174: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd192175: begin  
rid<=0;
end
19'd192301: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=65;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=22756;
 end   
19'd192302: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=55;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd192303: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=24;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd192304: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=93;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd192305: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=45;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd192306: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=24;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd192307: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=18;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd192308: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=85;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd192309: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=52;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd192310: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=98;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=39305;
 end   
19'd192311: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=70;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd192312: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=72;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd192313: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=66;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd192314: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=49;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd192315: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=59;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd192316: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=43;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd192317: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=85;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd192318: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=4;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd192319: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd192461: begin  
rid<=1;
end
19'd192462: begin  
end
19'd192463: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd192464: begin  
rid<=0;
end
19'd192601: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=31;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10675;
 end   
19'd192602: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=65;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd192603: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=79;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd192604: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=21;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd192605: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=11;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd192606: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=89;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=23680;
 end   
19'd192607: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=54;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd192608: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=17;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd192609: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=63;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd192610: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=53;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd192611: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd192753: begin  
rid<=1;
end
19'd192754: begin  
end
19'd192755: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd192756: begin  
rid<=0;
end
19'd192901: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=21;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=29235;
 end   
19'd192902: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=7;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=30900;
 end   
19'd192903: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=42;
   mapp<=39;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=23990;
 end   
19'd192904: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=58;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd192905: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=49;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd192906: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=96;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd192907: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=16;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd192908: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=49;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd192909: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=83;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd192910: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd192911: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd192912: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=84;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=51129;
 end   
19'd192913: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=60;
   mapp<=4;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=46981;
 end   
19'd192914: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=51;
   mapp<=42;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=46999;
 end   
19'd192915: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=64;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd192916: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=60;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd192917: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=84;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd192918: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=9;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd192919: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=68;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd192920: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=24;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd192921: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd192922: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd192923: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd193065: begin  
rid<=1;
end
19'd193066: begin  
end
19'd193067: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd193068: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd193069: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd193070: begin  
rid<=0;
end
19'd193201: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=92;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2300;
 end   
19'd193202: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=79;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7278;
 end   
19'd193203: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=67;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6184;
 end   
19'd193204: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=55;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5090;
 end   
19'd193205: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=57;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5284;
 end   
19'd193206: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=34;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=3178;
 end   
19'd193207: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=17;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=1624;
 end   
19'd193208: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=70;
 end   
19'd193209: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=40;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=3760;
 end   
19'd193210: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=23;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=2206;
 end   
19'd193211: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=53;
   pp<=100;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[10]<=4976;
 end   
19'd193212: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=18;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=2444;
 end   
19'd193213: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8286;
 end   
19'd193214: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=86;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=7732;
 end   
19'd193215: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=16;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=5378;
 end   
19'd193216: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=23;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=5698;
 end   
19'd193217: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=88;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=4762;
 end   
19'd193218: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=32;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=2200;
 end   
19'd193219: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=46;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=898;
 end   
19'd193220: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=74;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=5092;
 end   
19'd193221: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=61;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=3304;
 end   
19'd193222: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=23;
   pp<=100;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[10]<=5390;
 end   
19'd193223: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd193365: begin  
rid<=1;
end
19'd193366: begin  
end
19'd193367: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd193368: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd193369: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd193370: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd193371: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd193372: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd193373: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd193374: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd193375: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd193376: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd193377: begin  
check0<=expctdoutput[10]-outcheck0;
end
19'd193378: begin  
rid<=0;
end
19'd193501: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=33;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2211;
 end   
19'd193502: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=6;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=208;
 end   
19'd193503: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=55;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1835;
 end   
19'd193504: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=31;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1053;
 end   
19'd193505: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=80;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2680;
 end   
19'd193506: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=56;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=1898;
 end   
19'd193507: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=3;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=2460;
 end   
19'd193508: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=26;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=286;
 end   
19'd193509: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=74;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=2057;
 end   
19'd193510: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=89;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=1320;
 end   
19'd193511: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=46;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=2818;
 end   
19'd193512: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=65;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=2093;
 end   
19'd193513: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd193655: begin  
rid<=1;
end
19'd193656: begin  
end
19'd193657: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd193658: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd193659: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd193660: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd193661: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd193662: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd193663: begin  
rid<=0;
end
19'd193801: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=77;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9677;
 end   
19'd193802: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=87;
   mapp<=36;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4783;
 end   
19'd193803: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=23;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5793;
 end   
19'd193804: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=46;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4790;
 end   
19'd193805: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=14;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2597;
 end   
19'd193806: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=17;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=9276;
 end   
19'd193807: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=91;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=10373;
 end   
19'd193808: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=38;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=6998;
 end   
19'd193809: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=46;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=11713;
 end   
19'd193810: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=93;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=14733;
 end   
19'd193811: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd193812: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=33;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14984;
 end   
19'd193813: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=48;
   mapp<=81;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=9616;
 end   
19'd193814: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=45;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=8334;
 end   
19'd193815: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=22;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=9884;
 end   
19'd193816: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=91;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=7232;
 end   
19'd193817: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=34;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=14574;
 end   
19'd193818: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=87;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=17852;
 end   
19'd193819: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=96;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=13622;
 end   
19'd193820: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=72;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=17833;
 end   
19'd193821: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=78;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=19995;
 end   
19'd193822: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd193823: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd193965: begin  
rid<=1;
end
19'd193966: begin  
end
19'd193967: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd193968: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd193969: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd193970: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd193971: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd193972: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd193973: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd193974: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd193975: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd193976: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd193977: begin  
rid<=0;
end
19'd194101: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=14;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8831;
 end   
19'd194102: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=67;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8840;
 end   
19'd194103: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=40;
   mapp<=38;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8134;
 end   
19'd194104: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=28;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=12703;
 end   
19'd194105: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=81;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=15432;
 end   
19'd194106: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=84;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=13359;
 end   
19'd194107: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=67;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=9539;
 end   
19'd194108: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=51;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=4943;
 end   
19'd194109: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=17;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd194110: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=7;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd194111: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=27;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=15142;
 end   
19'd194112: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=68;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=16618;
 end   
19'd194113: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=22;
   mapp<=7;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15221;
 end   
19'd194114: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=90;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=21800;
 end   
19'd194115: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=19;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=19248;
 end   
19'd194116: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=29;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=20215;
 end   
19'd194117: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=77;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=16791;
 end   
19'd194118: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=3;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=8522;
 end   
19'd194119: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=55;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd194120: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd194121: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd194263: begin  
rid<=1;
end
19'd194264: begin  
end
19'd194265: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd194266: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd194267: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd194268: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd194269: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd194270: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd194271: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd194272: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd194273: begin  
rid<=0;
end
19'd194401: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=57;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12024;
 end   
19'd194402: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=90;
   mapp<=71;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11717;
 end   
19'd194403: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=25;
   mapp<=84;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7443;
 end   
19'd194404: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=4;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=9798;
 end   
19'd194405: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=91;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=12512;
 end   
19'd194406: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=54;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=14158;
 end   
19'd194407: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=97;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=14994;
 end   
19'd194408: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd194409: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd194410: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=27;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=25095;
 end   
19'd194411: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=78;
   mapp<=74;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=24207;
 end   
19'd194412: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=92;
   mapp<=72;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=21893;
 end   
19'd194413: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=53;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=24031;
 end   
19'd194414: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=91;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=25693;
 end   
19'd194415: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=62;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=26712;
 end   
19'd194416: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=64;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=27142;
 end   
19'd194417: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd194418: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd194419: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd194561: begin  
rid<=1;
end
19'd194562: begin  
end
19'd194563: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd194564: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd194565: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd194566: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd194567: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd194568: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd194569: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd194570: begin  
rid<=0;
end
19'd194701: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=63;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2520;
 end   
19'd194702: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=55;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2210;
 end   
19'd194703: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=38;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=3774;
 end   
19'd194704: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=36;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=3398;
 end   
19'd194705: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd194847: begin  
rid<=1;
end
19'd194848: begin  
end
19'd194849: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd194850: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd194851: begin  
rid<=0;
end
19'd195001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=46;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=414;
 end   
19'd195002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=75;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3460;
 end   
19'd195003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=41;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1906;
 end   
19'd195004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=78;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3618;
 end   
19'd195005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=56;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2616;
 end   
19'd195006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=62;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=2902;
 end   
19'd195007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=94;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=4384;
 end   
19'd195008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=57;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=2692;
 end   
19'd195009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=92;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=4312;
 end   
19'd195010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=52;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=2482;
 end   
19'd195011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=39;
   pp<=100;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[10]<=1894;
 end   
19'd195012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=51;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=3168;
 end   
19'd195013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=5092;
 end   
19'd195014: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=99;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=6955;
 end   
19'd195015: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=72;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=7290;
 end   
19'd195016: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=78;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=6594;
 end   
19'd195017: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=35;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=4687;
 end   
19'd195018: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=80;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=8464;
 end   
19'd195019: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=94;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=7486;
 end   
19'd195020: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=96;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=9208;
 end   
19'd195021: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=61;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=5593;
 end   
19'd195022: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=2;
   pp<=100;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[10]<=1996;
 end   
19'd195023: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd195165: begin  
rid<=1;
end
19'd195166: begin  
end
19'd195167: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd195168: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd195169: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd195170: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd195171: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd195172: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd195173: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd195174: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd195175: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd195176: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd195177: begin  
check0<=expctdoutput[10]-outcheck0;
end
19'd195178: begin  
rid<=0;
end
19'd195301: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=22;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11370;
 end   
19'd195302: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=5;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd195303: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd195304: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd195305: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=47;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd195306: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=57;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd195307: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=37;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd195308: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=77;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd195309: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=65;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=37993;
 end   
19'd195310: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=68;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd195311: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=97;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd195312: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=33;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd195313: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=91;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd195314: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=41;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd195315: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=21;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd195316: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=2;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd195317: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd195459: begin  
rid<=1;
end
19'd195460: begin  
end
19'd195461: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd195462: begin  
rid<=0;
end
19'd195601: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=38;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=888;
 end   
19'd195602: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=26;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=372;
 end   
19'd195603: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=11;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1218;
 end   
19'd195604: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=30;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1352;
 end   
19'd195605: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=7;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1060;
 end   
19'd195606: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=29;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=1152;
 end   
19'd195607: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=138;
 end   
19'd195608: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=3;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=1432;
 end   
19'd195609: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=48;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=1930;
 end   
19'd195610: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd195611: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=66;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=13524;
 end   
19'd195612: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=84;
   mapp<=86;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=9744;
 end   
19'd195613: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=44;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=11010;
 end   
19'd195614: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=82;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=8864;
 end   
19'd195615: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=25;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=9514;
 end   
19'd195616: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=81;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=6834;
 end   
19'd195617: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=4;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=1830;
 end   
19'd195618: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=17;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=10786;
 end   
19'd195619: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=98;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=11506;
 end   
19'd195620: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd195621: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd195763: begin  
rid<=1;
end
19'd195764: begin  
end
19'd195765: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd195766: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd195767: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd195768: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd195769: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd195770: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd195771: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd195772: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd195773: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd195774: begin  
rid<=0;
end
19'd195901: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=59;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=24160;
 end   
19'd195902: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=47;
   mapp<=86;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=25651;
 end   
19'd195903: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=62;
   mapp<=55;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=28515;
 end   
19'd195904: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=86;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd195905: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=62;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd195906: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=79;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd195907: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=83;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd195908: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=41;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd195909: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=2;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=33310;
 end   
19'd195910: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=53;
   mapp<=90;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=38501;
 end   
19'd195911: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=2;
   mapp<=22;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=39977;
 end   
19'd195912: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=8;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd195913: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=78;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd195914: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=69;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd195915: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=74;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd195916: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=80;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd195917: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd196059: begin  
rid<=1;
end
19'd196060: begin  
end
19'd196061: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd196062: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd196063: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd196064: begin  
rid<=0;
end
19'd196201: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=57;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=57;
 end   
19'd196202: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=93;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=103;
 end   
19'd196203: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=64;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=84;
 end   
19'd196204: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=69;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=99;
 end   
19'd196205: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=8;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=48;
 end   
19'd196206: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=77;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=127;
 end   
19'd196207: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=22;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=82;
 end   
19'd196208: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=97;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=167;
 end   
19'd196209: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=40;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=3497;
 end   
19'd196210: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=72;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=6295;
 end   
19'd196211: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=95;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=8254;
 end   
19'd196212: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=97;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=8441;
 end   
19'd196213: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=90;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=7788;
 end   
19'd196214: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=81;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=7093;
 end   
19'd196215: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=56;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=4898;
 end   
19'd196216: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=11;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=1113;
 end   
19'd196217: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd196359: begin  
rid<=1;
end
19'd196360: begin  
end
19'd196361: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd196362: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd196363: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd196364: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd196365: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd196366: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd196367: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd196368: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd196369: begin  
rid<=0;
end
19'd196501: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=6;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=996;
 end   
19'd196502: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=10;
   mapp<=78;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6532;
 end   
19'd196503: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=79;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10118;
 end   
19'd196504: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=93;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=11100;
 end   
19'd196505: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=99;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=10390;
 end   
19'd196506: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=87;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7784;
 end   
19'd196507: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=59;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=9516;
 end   
19'd196508: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=94;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=9850;
 end   
19'd196509: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=82;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd196510: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=0;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=1216;
 end   
19'd196511: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=10;
   mapp<=22;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=7600;
 end   
19'd196512: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=29;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=12553;
 end   
19'd196513: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=54;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=14368;
 end   
19'd196514: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=43;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=14197;
 end   
19'd196515: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=89;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=13239;
 end   
19'd196516: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=74;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=13490;
 end   
19'd196517: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=36;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=13114;
 end   
19'd196518: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=78;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd196519: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd196661: begin  
rid<=1;
end
19'd196662: begin  
end
19'd196663: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd196664: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd196665: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd196666: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd196667: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd196668: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd196669: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd196670: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd196671: begin  
rid<=0;
end
19'd196801: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=36;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13122;
 end   
19'd196802: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=3;
   mapp<=64;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=17788;
 end   
19'd196803: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=82;
   mapp<=53;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=19269;
 end   
19'd196804: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=80;
   mapp<=92;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=14102;
 end   
19'd196805: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=89;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=13794;
 end   
19'd196806: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=72;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=10465;
 end   
19'd196807: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=20;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=7077;
 end   
19'd196808: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=55;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=8891;
 end   
19'd196809: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=41;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd196810: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=7;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd196811: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=43;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd196812: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=49;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=19958;
 end   
19'd196813: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=31;
   mapp<=21;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=29364;
 end   
19'd196814: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=99;
   mapp<=34;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=27784;
 end   
19'd196815: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=12;
   mapp<=92;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=25769;
 end   
19'd196816: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=87;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=28217;
 end   
19'd196817: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=20;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=18132;
 end   
19'd196818: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=95;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=13960;
 end   
19'd196819: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=84;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=16368;
 end   
19'd196820: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd196821: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=11;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd196822: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=40;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd196823: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd196965: begin  
rid<=1;
end
19'd196966: begin  
end
19'd196967: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd196968: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd196969: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd196970: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd196971: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd196972: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd196973: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd196974: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd196975: begin  
rid<=0;
end
19'd197101: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=71;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7722;
 end   
19'd197102: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=67;
   mapp<=79;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8981;
 end   
19'd197103: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=90;
   mapp<=12;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5649;
 end   
19'd197104: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=49;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1289;
 end   
19'd197105: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=4;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1107;
 end   
19'd197106: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=1;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7093;
 end   
19'd197107: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=76;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=9299;
 end   
19'd197108: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=85;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=8891;
 end   
19'd197109: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=90;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=2974;
 end   
19'd197110: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=8;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd197111: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=46;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd197112: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=32;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=11096;
 end   
19'd197113: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=42;
   mapp<=61;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12471;
 end   
19'd197114: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=26;
   mapp<=14;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=11873;
 end   
19'd197115: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=94;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=3924;
 end   
19'd197116: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=9;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=5890;
 end   
19'd197117: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=55;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=14390;
 end   
19'd197118: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=93;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=14770;
 end   
19'd197119: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=61;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=11809;
 end   
19'd197120: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=32;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=4204;
 end   
19'd197121: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=8;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd197122: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=21;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd197123: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd197265: begin  
rid<=1;
end
19'd197266: begin  
end
19'd197267: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd197268: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd197269: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd197270: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd197271: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd197272: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd197273: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd197274: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd197275: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd197276: begin  
rid<=0;
end
19'd197401: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=24;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7645;
 end   
19'd197402: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=12;
   mapp<=33;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8068;
 end   
19'd197403: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=49;
   mapp<=81;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5975;
 end   
19'd197404: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=61;
   mapp<=40;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4297;
 end   
19'd197405: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=27;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5127;
 end   
19'd197406: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=1;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=5406;
 end   
19'd197407: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=29;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd197408: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=44;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd197409: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=20;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd197410: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=25;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14107;
 end   
19'd197411: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=44;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=14554;
 end   
19'd197412: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=62;
   mapp<=32;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15194;
 end   
19'd197413: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=9;
   mapp<=77;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=9985;
 end   
19'd197414: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=2;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=15709;
 end   
19'd197415: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=49;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=17581;
 end   
19'd197416: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=43;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd197417: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=92;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd197418: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=46;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd197419: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd197561: begin  
rid<=1;
end
19'd197562: begin  
end
19'd197563: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd197564: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd197565: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd197566: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd197567: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd197568: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd197569: begin  
rid<=0;
end
19'd197701: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=48;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3527;
 end   
19'd197702: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=5;
   mapp<=16;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2415;
 end   
19'd197703: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=23;
   mapp<=33;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3258;
 end   
19'd197704: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd197705: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd197706: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=62;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12938;
 end   
19'd197707: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=81;
   mapp<=81;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=15907;
 end   
19'd197708: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=76;
   mapp<=22;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=12738;
 end   
19'd197709: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd197710: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd197711: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd197853: begin  
rid<=1;
end
19'd197854: begin  
end
19'd197855: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd197856: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd197857: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd197858: begin  
rid<=0;
end
19'd198001: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=72;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=31003;
 end   
19'd198002: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=71;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd198003: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=4;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd198004: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=91;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd198005: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=82;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd198006: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=93;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd198007: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=24;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd198008: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=67;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd198009: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=47;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd198010: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=67;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=60225;
 end   
19'd198011: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=53;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd198012: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=77;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd198013: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=1;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd198014: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=95;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd198015: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=38;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd198016: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=35;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd198017: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=85;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd198018: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=91;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd198019: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd198161: begin  
rid<=1;
end
19'd198162: begin  
end
19'd198163: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd198164: begin  
rid<=0;
end
19'd198301: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=62;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10549;
 end   
19'd198302: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=30;
   mapp<=96;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11040;
 end   
19'd198303: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=4;
   mapp<=97;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12494;
 end   
19'd198304: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=73;
   mapp<=25;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=17873;
 end   
19'd198305: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=37;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=18593;
 end   
19'd198306: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=61;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=21756;
 end   
19'd198307: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=78;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd198308: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=75;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd198309: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=63;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd198310: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=71;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=21508;
 end   
19'd198311: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=43;
   mapp<=99;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=24922;
 end   
19'd198312: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=98;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=35108;
 end   
19'd198313: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=82;
   mapp<=80;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=38919;
 end   
19'd198314: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=72;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=36988;
 end   
19'd198315: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=93;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=32920;
 end   
19'd198316: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=58;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd198317: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=42;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd198318: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=14;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd198319: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd198461: begin  
rid<=1;
end
19'd198462: begin  
end
19'd198463: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd198464: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd198465: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd198466: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd198467: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd198468: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd198469: begin  
rid<=0;
end
19'd198601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=54;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12485;
 end   
19'd198602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=71;
   mapp<=29;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12065;
 end   
19'd198603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=76;
   mapp<=91;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=14397;
 end   
19'd198604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=53;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=10725;
 end   
19'd198605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=75;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=7649;
 end   
19'd198606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd198607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd198608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=94;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=21855;
 end   
19'd198609: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=69;
   mapp<=71;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=24829;
 end   
19'd198610: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=9;
   mapp<=79;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=27199;
 end   
19'd198611: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=71;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=21821;
 end   
19'd198612: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=53;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=18901;
 end   
19'd198613: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd198614: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd198615: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd198757: begin  
rid<=1;
end
19'd198758: begin  
end
19'd198759: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd198760: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd198761: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd198762: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd198763: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd198764: begin  
rid<=0;
end
19'd198901: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=77;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5339;
 end   
19'd198902: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=15;
   mapp<=89;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7958;
 end   
19'd198903: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=73;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6436;
 end   
19'd198904: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=53;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4651;
 end   
19'd198905: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd198906: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=10907;
 end   
19'd198907: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=64;
   mapp<=87;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=11542;
 end   
19'd198908: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=56;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=7588;
 end   
19'd198909: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=18;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=5227;
 end   
19'd198910: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd198911: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd199053: begin  
rid<=1;
end
19'd199054: begin  
end
19'd199055: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd199056: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd199057: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd199058: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd199059: begin  
rid<=0;
end
19'd199201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=74;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9253;
 end   
19'd199202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=97;
   mapp<=66;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8709;
 end   
19'd199203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=83;
   mapp<=29;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6611;
 end   
19'd199204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=91;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd199205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=3;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd199206: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=32;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=20204;
 end   
19'd199207: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=97;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=19397;
 end   
19'd199208: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=51;
   mapp<=69;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=16679;
 end   
19'd199209: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=82;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd199210: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=50;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd199211: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd199353: begin  
rid<=1;
end
19'd199354: begin  
end
19'd199355: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd199356: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd199357: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd199358: begin  
rid<=0;
end
19'd199501: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=74;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=27908;
 end   
19'd199502: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=28;
   mapp<=66;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=25481;
 end   
19'd199503: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=17;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd199504: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=86;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd199505: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=62;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd199506: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=29;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd199507: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=72;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd199508: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=89;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd199509: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=91;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd199510: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=22;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd199511: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd199512: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=86;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=70385;
 end   
19'd199513: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=83;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=72278;
 end   
19'd199514: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=71;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd199515: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=98;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd199516: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=94;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd199517: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=69;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd199518: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=59;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd199519: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=84;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd199520: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=48;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd199521: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=68;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd199522: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd199523: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd199665: begin  
rid<=1;
end
19'd199666: begin  
end
19'd199667: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd199668: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd199669: begin  
rid<=0;
end
19'd199801: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=89;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=17423;
 end   
19'd199802: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=7;
   mapp<=43;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=23005;
 end   
19'd199803: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=61;
   mapp<=81;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=27193;
 end   
19'd199804: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=55;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd199805: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=41;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd199806: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=14;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd199807: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=94;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd199808: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=77;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd199809: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd199810: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd199811: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=90;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=47091;
 end   
19'd199812: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=7;
   mapp<=82;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=55494;
 end   
19'd199813: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=88;
   mapp<=16;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=51885;
 end   
19'd199814: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=58;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd199815: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=53;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd199816: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=45;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd199817: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=83;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd199818: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=92;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd199819: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd199820: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd199821: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd199963: begin  
rid<=1;
end
19'd199964: begin  
end
19'd199965: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd199966: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd199967: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd199968: begin  
rid<=0;
end
19'd200101: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=43;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10468;
 end   
19'd200102: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=17;
   mapp<=16;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12385;
 end   
19'd200103: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=62;
   mapp<=94;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11122;
 end   
19'd200104: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=4;
   mapp<=91;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=10289;
 end   
19'd200105: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=65;
   mapp<=28;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6991;
 end   
19'd200106: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd200107: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=15;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd200108: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd200109: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd200110: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd200111: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd200112: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=78;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=24476;
 end   
19'd200113: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=15;
   mapp<=8;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=22154;
 end   
19'd200114: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=11;
   mapp<=75;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=25410;
 end   
19'd200115: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=80;
   mapp<=86;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=26566;
 end   
19'd200116: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=34;
   mapp<=27;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=17768;
 end   
19'd200117: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=24;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd200118: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=39;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd200119: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd200120: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd200121: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd200122: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd200123: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd200265: begin  
rid<=1;
end
19'd200266: begin  
end
19'd200267: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd200268: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd200269: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd200270: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd200271: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd200272: begin  
rid<=0;
end
19'd200401: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=11;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=15018;
 end   
19'd200402: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=59;
   mapp<=6;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=21823;
 end   
19'd200403: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=83;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd200404: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=85;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd200405: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=2;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd200406: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=89;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd200407: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=48;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd200408: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=2;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd200409: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=64;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd200410: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd200411: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=20;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=30387;
 end   
19'd200412: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=16;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=37054;
 end   
19'd200413: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=36;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd200414: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=95;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd200415: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=39;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd200416: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=74;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd200417: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=22;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd200418: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=17;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd200419: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=16;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd200420: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd200421: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd200563: begin  
rid<=1;
end
19'd200564: begin  
end
19'd200565: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd200566: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd200567: begin  
rid<=0;
end
19'd200701: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=69;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4257;
 end   
19'd200702: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=31;
   mapp<=92;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9963;
 end   
19'd200703: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=38;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd200704: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd200705: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=95;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=27139;
 end   
19'd200706: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=98;
   mapp<=96;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=32711;
 end   
19'd200707: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=68;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd200708: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd200709: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd200851: begin  
rid<=1;
end
19'd200852: begin  
end
19'd200853: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd200854: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd200855: begin  
rid<=0;
end
19'd201001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=19;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4531;
 end   
19'd201002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=36;
   mapp<=28;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6922;
 end   
19'd201003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=28;
   mapp<=95;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7754;
 end   
19'd201004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=3;
   mapp<=95;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=2674;
 end   
19'd201005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=54;
   mapp<=10;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3892;
 end   
19'd201006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=5;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=3914;
 end   
19'd201007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=41;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=2301;
 end   
19'd201008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd201009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd201010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd201011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd201012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=8;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=19378;
 end   
19'd201013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=28;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=16295;
 end   
19'd201014: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=66;
   mapp<=91;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15275;
 end   
19'd201015: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=10;
   mapp<=79;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=7382;
 end   
19'd201016: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=75;
   mapp<=61;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=11131;
 end   
19'd201017: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=3;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=9547;
 end   
19'd201018: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=7;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=13450;
 end   
19'd201019: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd201020: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd201021: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd201022: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd201023: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd201165: begin  
rid<=1;
end
19'd201166: begin  
end
19'd201167: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd201168: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd201169: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd201170: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd201171: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd201172: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd201173: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd201174: begin  
rid<=0;
end
19'd201301: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=59;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7730;
 end   
19'd201302: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=68;
   mapp<=46;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7844;
 end   
19'd201303: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=55;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd201304: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=78;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=15213;
 end   
19'd201305: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=77;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=15811;
 end   
19'd201306: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=83;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd201307: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd201449: begin  
rid<=1;
end
19'd201450: begin  
end
19'd201451: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd201452: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd201453: begin  
rid<=0;
end
19'd201601: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=4;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13322;
 end   
19'd201602: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=88;
   mapp<=96;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7339;
 end   
19'd201603: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=69;
   mapp<=68;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2609;
 end   
19'd201604: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=26;
   mapp<=3;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3148;
 end   
19'd201605: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=29;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1930;
 end   
19'd201606: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd201607: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd201608: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd201609: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=85;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=21188;
 end   
19'd201610: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=30;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=14143;
 end   
19'd201611: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=21;
   mapp<=51;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=10570;
 end   
19'd201612: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=80;
   mapp<=34;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=8949;
 end   
19'd201613: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=6;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=8156;
 end   
19'd201614: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd201615: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd201616: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd201617: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd201759: begin  
rid<=1;
end
19'd201760: begin  
end
19'd201761: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd201762: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd201763: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd201764: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd201765: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd201766: begin  
rid<=0;
end
19'd201901: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=43;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2734;
 end   
19'd201902: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=33;
   mapp<=17;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1509;
 end   
19'd201903: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=1;
   mapp<=23;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1329;
 end   
19'd201904: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=9;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1195;
 end   
19'd201905: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=23;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1672;
 end   
19'd201906: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=19;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=1428;
 end   
19'd201907: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=16;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=1871;
 end   
19'd201908: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=33;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=2636;
 end   
19'd201909: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd201910: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd201911: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=99;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12230;
 end   
19'd201912: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=51;
   mapp<=26;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=10538;
 end   
19'd201913: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=47;
   mapp<=98;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=16231;
 end   
19'd201914: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=31;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=9366;
 end   
19'd201915: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=77;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=11275;
 end   
19'd201916: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=25;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=5890;
 end   
19'd201917: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=15;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=8724;
 end   
19'd201918: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=26;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=10959;
 end   
19'd201919: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd201920: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd201921: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd202063: begin  
rid<=1;
end
19'd202064: begin  
end
19'd202065: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd202066: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd202067: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd202068: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd202069: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd202070: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd202071: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd202072: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd202073: begin  
rid<=0;
end
19'd202201: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=9;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=387;
 end   
19'd202202: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=2;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=96;
 end   
19'd202203: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=91;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3933;
 end   
19'd202204: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=73;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3169;
 end   
19'd202205: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=94;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4082;
 end   
19'd202206: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=79;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=3447;
 end   
19'd202207: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=2;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=146;
 end   
19'd202208: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=75;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=3295;
 end   
19'd202209: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=86;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5891;
 end   
19'd202210: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=86;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=5600;
 end   
19'd202211: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=90;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=9693;
 end   
19'd202212: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=58;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6881;
 end   
19'd202213: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=65;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=8242;
 end   
19'd202214: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=3447;
 end   
19'd202215: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=64;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=4242;
 end   
19'd202216: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=71;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=7839;
 end   
19'd202217: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd202359: begin  
rid<=1;
end
19'd202360: begin  
end
19'd202361: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd202362: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd202363: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd202364: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd202365: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd202366: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd202367: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd202368: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd202369: begin  
rid<=0;
end
19'd202501: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=93;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8277;
 end   
19'd202502: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=0;
   mapp<=70;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6520;
 end   
19'd202503: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=5;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8517;
 end   
19'd202504: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=0;
   mapp<=21;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=6625;
 end   
19'd202505: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd202647: begin  
rid<=1;
end
19'd202648: begin  
end
19'd202649: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd202650: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd202651: begin  
rid<=0;
end
19'd202801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=2;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8666;
 end   
19'd202802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=7;
   mapp<=42;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2927;
 end   
19'd202803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=97;
   mapp<=86;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=935;
 end   
19'd202804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=23;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=8945;
 end   
19'd202805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=6;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=7479;
 end   
19'd202806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd202807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd202808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=84;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12406;
 end   
19'd202809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=14;
   mapp<=74;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=11038;
 end   
19'd202810: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=37;
   mapp<=64;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=8539;
 end   
19'd202811: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=27;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=14392;
 end   
19'd202812: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=50;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=13764;
 end   
19'd202813: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd202814: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd202815: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd202957: begin  
rid<=1;
end
19'd202958: begin  
end
19'd202959: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd202960: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd202961: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd202962: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd202963: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd202964: begin  
rid<=0;
end
19'd203101: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=69;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8188;
 end   
19'd203102: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=6;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=13606;
 end   
19'd203103: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=64;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd203104: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd203105: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=55;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=15798;
 end   
19'd203106: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=9;
   mapp<=15;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20842;
 end   
19'd203107: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=85;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd203108: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=69;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd203109: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd203251: begin  
rid<=1;
end
19'd203252: begin  
end
19'd203253: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd203254: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd203255: begin  
rid<=0;
end
19'd203401: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=9;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=288;
 end   
19'd203402: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=75;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=685;
 end   
19'd203403: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=4;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=56;
 end   
19'd203404: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=30;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=300;
 end   
19'd203405: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=80;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=760;
 end   
19'd203406: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=7;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=113;
 end   
19'd203407: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=92;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=888;
 end   
19'd203408: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=90;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=880;
 end   
19'd203409: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=28;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=332;
 end   
19'd203410: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=75;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=765;
 end   
19'd203411: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=82;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8324;
 end   
19'd203412: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=31;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=3227;
 end   
19'd203413: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=82;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=6780;
 end   
19'd203414: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=30;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=2760;
 end   
19'd203415: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=35;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=3630;
 end   
19'd203416: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=6;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=605;
 end   
19'd203417: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=64;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=6136;
 end   
19'd203418: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=5;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=1290;
 end   
19'd203419: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=18;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=1808;
 end   
19'd203420: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=22;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=2569;
 end   
19'd203421: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd203563: begin  
rid<=1;
end
19'd203564: begin  
end
19'd203565: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd203566: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd203567: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd203568: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd203569: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd203570: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd203571: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd203572: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd203573: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd203574: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd203575: begin  
rid<=0;
end
19'd203701: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=78;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8717;
 end   
19'd203702: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=25;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6241;
 end   
19'd203703: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=44;
   mapp<=9;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4550;
 end   
19'd203704: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5681;
 end   
19'd203705: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=87;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=9857;
 end   
19'd203706: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=79;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=10420;
 end   
19'd203707: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd203708: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd203709: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=75;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14104;
 end   
19'd203710: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=8;
   mapp<=73;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12399;
 end   
19'd203711: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=51;
   mapp<=28;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=9986;
 end   
19'd203712: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=9;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=10846;
 end   
19'd203713: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=64;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=18902;
 end   
19'd203714: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=78;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=18929;
 end   
19'd203715: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd203716: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd203717: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd203859: begin  
rid<=1;
end
19'd203860: begin  
end
19'd203861: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd203862: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd203863: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd203864: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd203865: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd203866: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd203867: begin  
rid<=0;
end
19'd204001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=99;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9172;
 end   
19'd204002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=80;
   mapp<=31;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8381;
 end   
19'd204003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=21;
   mapp<=24;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10470;
 end   
19'd204004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=20;
   mapp<=45;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=12367;
 end   
19'd204005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=16;
   mapp<=83;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=12167;
 end   
19'd204006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=40;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=9231;
 end   
19'd204007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=82;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=9343;
 end   
19'd204008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=77;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd204009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=58;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd204010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=7;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd204011: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd204012: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=3;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17461;
 end   
19'd204013: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=43;
   mapp<=24;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=19460;
 end   
19'd204014: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=24;
   mapp<=68;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=22070;
 end   
19'd204015: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=55;
   mapp<=78;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=26692;
 end   
19'd204016: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=34;
   mapp<=36;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=25143;
 end   
19'd204017: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=70;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=20795;
 end   
19'd204018: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=45;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=17430;
 end   
19'd204019: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd204020: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=1;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd204021: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=49;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd204022: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=11;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd204023: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd204165: begin  
rid<=1;
end
19'd204166: begin  
end
19'd204167: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd204168: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd204169: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd204170: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd204171: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd204172: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd204173: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd204174: begin  
rid<=0;
end
19'd204301: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=96;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=17401;
 end   
19'd204302: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=53;
   mapp<=58;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10742;
 end   
19'd204303: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=50;
   mapp<=18;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7457;
 end   
19'd204304: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=5;
   mapp<=18;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=9003;
 end   
19'd204305: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=77;
   mapp<=61;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=10495;
 end   
19'd204306: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=26;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=4917;
 end   
19'd204307: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=13;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=9086;
 end   
19'd204308: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=55;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd204309: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=13;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd204310: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=9;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd204311: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd204312: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=84;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=38240;
 end   
19'd204313: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=54;
   mapp<=81;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=24252;
 end   
19'd204314: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=41;
   mapp<=41;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=22889;
 end   
19'd204315: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=36;
   mapp<=5;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=23275;
 end   
19'd204316: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=83;
   mapp<=96;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=25221;
 end   
19'd204317: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=42;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=15141;
 end   
19'd204318: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=59;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=20459;
 end   
19'd204319: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=28;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd204320: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd204321: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=9;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd204322: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=36;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd204323: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd204465: begin  
rid<=1;
end
19'd204466: begin  
end
19'd204467: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd204468: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd204469: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd204470: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd204471: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd204472: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd204473: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd204474: begin  
rid<=0;
end
19'd204601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=48;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=17558;
 end   
19'd204602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=28;
   mapp<=16;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=21976;
 end   
19'd204603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=61;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd204604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=46;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd204605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=85;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd204606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=93;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd204607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd204608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=76;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=36873;
 end   
19'd204609: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=87;
   mapp<=42;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=39443;
 end   
19'd204610: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=71;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd204611: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=45;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd204612: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=14;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd204613: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=31;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd204614: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd204615: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd204757: begin  
rid<=1;
end
19'd204758: begin  
end
19'd204759: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd204760: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd204761: begin  
rid<=0;
end
19'd204901: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=99;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4851;
 end   
19'd204902: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4762;
 end   
19'd204903: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=97;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9623;
 end   
19'd204904: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=62;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6168;
 end   
19'd204905: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=62;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6178;
 end   
19'd204906: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=44;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=4406;
 end   
19'd204907: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=95;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=9465;
 end   
19'd204908: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=91;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=9079;
 end   
19'd204909: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=68;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7027;
 end   
19'd204910: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=78;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=10066;
 end   
19'd204911: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=79;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=14995;
 end   
19'd204912: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=93;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=12492;
 end   
19'd204913: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=25;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=7878;
 end   
19'd204914: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=32;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=6582;
 end   
19'd204915: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=33;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=11709;
 end   
19'd204916: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=95;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=15539;
 end   
19'd204917: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd205059: begin  
rid<=1;
end
19'd205060: begin  
end
19'd205061: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd205062: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd205063: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd205064: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd205065: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd205066: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd205067: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd205068: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd205069: begin  
rid<=0;
end
19'd205201: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=58;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=28718;
 end   
19'd205202: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=68;
   mapp<=52;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=20204;
 end   
19'd205203: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=94;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd205204: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=10;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd205205: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=90;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd205206: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=54;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd205207: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=18;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd205208: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=62;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd205209: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=28;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd205210: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=68;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd205211: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=57;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=49195;
 end   
19'd205212: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=2;
   mapp<=13;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=34508;
 end   
19'd205213: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=13;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd205214: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=7;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd205215: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=71;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd205216: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=81;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd205217: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=3;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd205218: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=38;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd205219: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=24;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd205220: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd205221: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd205363: begin  
rid<=1;
end
19'd205364: begin  
end
19'd205365: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd205366: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd205367: begin  
rid<=0;
end
19'd205501: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=55;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=15453;
 end   
19'd205502: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=20;
   mapp<=26;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10087;
 end   
19'd205503: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=97;
   mapp<=94;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=14537;
 end   
19'd205504: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=38;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd205505: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=11;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd205506: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd205507: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd205508: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=65;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=28265;
 end   
19'd205509: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=88;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20743;
 end   
19'd205510: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=6;
   mapp<=20;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=25046;
 end   
19'd205511: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=25;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd205512: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=3;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd205513: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd205514: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd205515: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd205657: begin  
rid<=1;
end
19'd205658: begin  
end
19'd205659: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd205660: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd205661: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd205662: begin  
rid<=0;
end
19'd205801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=27;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=19443;
 end   
19'd205802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=30;
   mapp<=70;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=25887;
 end   
19'd205803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=65;
   mapp<=31;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=26855;
 end   
19'd205804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=70;
   mapp<=59;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=29605;
 end   
19'd205805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=71;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd205806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=32;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd205807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=95;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd205808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=64;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd205809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=93;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd205810: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=44;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd205811: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=78;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=33927;
 end   
19'd205812: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=37;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=39317;
 end   
19'd205813: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=4;
   mapp<=73;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=42247;
 end   
19'd205814: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=31;
   mapp<=11;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=45031;
 end   
19'd205815: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=57;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd205816: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=56;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd205817: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=73;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd205818: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=63;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd205819: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=53;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd205820: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=1;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd205821: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd205963: begin  
rid<=1;
end
19'd205964: begin  
end
19'd205965: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd205966: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd205967: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd205968: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd205969: begin  
rid<=0;
end
19'd206101: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=86;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3854;
 end   
19'd206102: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=93;
   mapp<=10;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3222;
 end   
19'd206103: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=5;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=610;
 end   
19'd206104: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=42;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd206105: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=39;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=10796;
 end   
19'd206106: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=40;
   mapp<=78;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=10418;
 end   
19'd206107: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=42;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=12214;
 end   
19'd206108: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=96;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd206109: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd206251: begin  
rid<=1;
end
19'd206252: begin  
end
19'd206253: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd206254: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd206255: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd206256: begin  
rid<=0;
end
19'd206401: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=17;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=629;
 end   
19'd206402: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=8;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=306;
 end   
19'd206403: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=24;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=908;
 end   
19'd206404: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=45;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1695;
 end   
19'd206405: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=80;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3000;
 end   
19'd206406: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=16;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=642;
 end   
19'd206407: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=89;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=3353;
 end   
19'd206408: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=49;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=1658;
 end   
19'd206409: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=16;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=642;
 end   
19'd206410: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=44;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=1832;
 end   
19'd206411: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=37;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=2472;
 end   
19'd206412: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=8;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=3168;
 end   
19'd206413: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=44;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=1566;
 end   
19'd206414: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=35;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=4088;
 end   
19'd206415: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd206557: begin  
rid<=1;
end
19'd206558: begin  
end
19'd206559: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd206560: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd206561: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd206562: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd206563: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd206564: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd206565: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd206566: begin  
rid<=0;
end
19'd206701: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=93;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14898;
 end   
19'd206702: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=9;
   mapp<=8;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8448;
 end   
19'd206703: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=16;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9366;
 end   
19'd206704: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=58;
   mapp<=62;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7624;
 end   
19'd206705: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=71;
   mapp<=90;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=15094;
 end   
19'd206706: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=12;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7068;
 end   
19'd206707: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=2;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=8766;
 end   
19'd206708: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd206709: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd206710: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd206711: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd206712: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=32;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=29254;
 end   
19'd206713: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=80;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=23343;
 end   
19'd206714: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=8;
   mapp<=93;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=25063;
 end   
19'd206715: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=79;
   mapp<=72;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=18506;
 end   
19'd206716: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=52;
   mapp<=29;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=25653;
 end   
19'd206717: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=47;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=19926;
 end   
19'd206718: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=58;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=15489;
 end   
19'd206719: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd206720: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd206721: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd206722: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd206723: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd206865: begin  
rid<=1;
end
19'd206866: begin  
end
19'd206867: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd206868: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd206869: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd206870: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd206871: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd206872: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd206873: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd206874: begin  
rid<=0;
end
19'd207001: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=69;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1344;
 end   
19'd207002: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=15;
   mapp<=85;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7760;
 end   
19'd207003: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=91;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6911;
 end   
19'd207004: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=80;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd207005: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=60;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5649;
 end   
19'd207006: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=45;
   mapp<=9;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=11036;
 end   
19'd207007: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=39;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=10274;
 end   
19'd207008: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=92;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd207009: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd207151: begin  
rid<=1;
end
19'd207152: begin  
end
19'd207153: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd207154: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd207155: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd207156: begin  
rid<=0;
end
19'd207301: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=66;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=21530;
 end   
19'd207302: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=88;
   mapp<=91;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=18186;
 end   
19'd207303: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=88;
   mapp<=58;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=18501;
 end   
19'd207304: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=61;
   mapp<=7;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=21294;
 end   
19'd207305: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=7;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd207306: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=68;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd207307: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=73;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd207308: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=4;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd207309: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd207310: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd207311: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd207312: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=55;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=41700;
 end   
19'd207313: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=16;
   mapp<=38;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=37960;
 end   
19'd207314: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=61;
   mapp<=23;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=41422;
 end   
19'd207315: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=54;
   mapp<=36;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=44789;
 end   
19'd207316: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=54;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd207317: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=96;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd207318: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=38;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd207319: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=1;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd207320: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd207321: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd207322: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd207323: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd207465: begin  
rid<=1;
end
19'd207466: begin  
end
19'd207467: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd207468: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd207469: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd207470: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd207471: begin  
rid<=0;
end
19'd207601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=42;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=22445;
 end   
19'd207602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=78;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd207603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=56;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd207604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=87;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd207605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=76;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd207606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=38;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd207607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=77;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd207608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=96;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=55621;
 end   
19'd207609: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=80;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd207610: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=82;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd207611: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=46;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd207612: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=98;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd207613: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=18;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd207614: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=85;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd207615: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd207757: begin  
rid<=1;
end
19'd207758: begin  
end
19'd207759: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd207760: begin  
rid<=0;
end
19'd207901: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=3;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=57;
 end   
19'd207902: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=85;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1625;
 end   
19'd207903: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=75;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1445;
 end   
19'd207904: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=58;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=3885;
 end   
19'd207905: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=69;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=6179;
 end   
19'd207906: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=6;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=1841;
 end   
19'd207907: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd208049: begin  
rid<=1;
end
19'd208050: begin  
end
19'd208051: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd208052: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd208053: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd208054: begin  
rid<=0;
end
19'd208201: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=55;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6290;
 end   
19'd208202: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=24;
   mapp<=18;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7072;
 end   
19'd208203: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=54;
   mapp<=82;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7434;
 end   
19'd208204: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=76;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=8740;
 end   
19'd208205: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=20;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5640;
 end   
19'd208206: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=75;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=8561;
 end   
19'd208207: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=50;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=6602;
 end   
19'd208208: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=59;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=4749;
 end   
19'd208209: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd208210: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd208211: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=97;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=15707;
 end   
19'd208212: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=24;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=17724;
 end   
19'd208213: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=48;
   mapp<=47;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=17201;
 end   
19'd208214: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=61;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=20033;
 end   
19'd208215: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=78;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=19662;
 end   
19'd208216: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=73;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=20874;
 end   
19'd208217: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=98;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=20812;
 end   
19'd208218: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=60;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=15849;
 end   
19'd208219: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd208220: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd208221: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd208363: begin  
rid<=1;
end
19'd208364: begin  
end
19'd208365: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd208366: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd208367: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd208368: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd208369: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd208370: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd208371: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd208372: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd208373: begin  
rid<=0;
end
19'd208501: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=77;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4466;
 end   
19'd208502: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=75;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5785;
 end   
19'd208503: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=67;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5179;
 end   
19'd208504: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=90;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6960;
 end   
19'd208505: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=58;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4506;
 end   
19'd208506: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=47;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=4701;
 end   
19'd208507: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=20;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=6725;
 end   
19'd208508: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=12;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=5743;
 end   
19'd208509: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=91;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=11237;
 end   
19'd208510: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=50;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=6856;
 end   
19'd208511: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd208653: begin  
rid<=1;
end
19'd208654: begin  
end
19'd208655: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd208656: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd208657: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd208658: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd208659: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd208660: begin  
rid<=0;
end
19'd208801: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=19;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9341;
 end   
19'd208802: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=44;
   mapp<=90;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12365;
 end   
19'd208803: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=34;
   mapp<=50;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10744;
 end   
19'd208804: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=33;
   mapp<=77;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=15081;
 end   
19'd208805: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=65;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=13473;
 end   
19'd208806: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=32;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=15880;
 end   
19'd208807: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=73;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=18919;
 end   
19'd208808: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=39;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd208809: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd208810: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=97;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd208811: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=56;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16997;
 end   
19'd208812: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=48;
   mapp<=52;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=19813;
 end   
19'd208813: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=64;
   mapp<=34;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=18096;
 end   
19'd208814: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=36;
   mapp<=16;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=21741;
 end   
19'd208815: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=52;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=20091;
 end   
19'd208816: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=60;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=22132;
 end   
19'd208817: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=23;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=24930;
 end   
19'd208818: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=30;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd208819: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=91;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd208820: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd208821: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd208963: begin  
rid<=1;
end
19'd208964: begin  
end
19'd208965: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd208966: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd208967: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd208968: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd208969: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd208970: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd208971: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd208972: begin  
rid<=0;
end
19'd209101: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=52;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14644;
 end   
19'd209102: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=91;
   mapp<=29;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12770;
 end   
19'd209103: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=27;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=17754;
 end   
19'd209104: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=35;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd209105: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=72;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd209106: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=74;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd209107: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=73;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd209108: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=6;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd209109: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd209110: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd209111: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=8;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=40883;
 end   
19'd209112: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=73;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=34843;
 end   
19'd209113: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=9;
   mapp<=49;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=44306;
 end   
19'd209114: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=72;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd209115: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=25;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd209116: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=87;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd209117: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=91;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd209118: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=42;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd209119: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd209120: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd209121: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd209263: begin  
rid<=1;
end
19'd209264: begin  
end
19'd209265: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd209266: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd209267: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd209268: begin  
rid<=0;
end
19'd209401: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=33;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9708;
 end   
19'd209402: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=8;
   mapp<=12;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10082;
 end   
19'd209403: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=59;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd209404: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=97;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd209405: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=79;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd209406: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd209407: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=57;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=20960;
 end   
19'd209408: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=4;
   mapp<=49;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18864;
 end   
19'd209409: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=65;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd209410: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=59;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd209411: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=6;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd209412: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd209413: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd209555: begin  
rid<=1;
end
19'd209556: begin  
end
19'd209557: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd209558: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd209559: begin  
rid<=0;
end
19'd209701: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=83;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5677;
 end   
19'd209702: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=49;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11267;
 end   
19'd209703: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=12;
   mapp<=93;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6317;
 end   
19'd209704: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=93;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=11005;
 end   
19'd209705: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=56;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=9498;
 end   
19'd209706: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=63;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=10171;
 end   
19'd209707: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=67;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=9939;
 end   
19'd209708: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd209709: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=65;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd209710: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=39;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=18062;
 end   
19'd209711: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=75;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=25811;
 end   
19'd209712: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=86;
   mapp<=44;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=18348;
 end   
19'd209713: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=83;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=19895;
 end   
19'd209714: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=24;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=19659;
 end   
19'd209715: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=85;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=19578;
 end   
19'd209716: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=25;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=20338;
 end   
19'd209717: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=93;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd209718: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd209719: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd209861: begin  
rid<=1;
end
19'd209862: begin  
end
19'd209863: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd209864: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd209865: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd209866: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd209867: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd209868: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd209869: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd209870: begin  
rid<=0;
end
19'd210001: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=84;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=20650;
 end   
19'd210002: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=45;
   mapp<=24;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=19541;
 end   
19'd210003: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=45;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd210004: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=24;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd210005: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=94;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd210006: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=4;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd210007: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=33;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd210008: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd210009: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=20;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=40201;
 end   
19'd210010: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=8;
   mapp<=24;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=33814;
 end   
19'd210011: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=41;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd210012: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=19;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd210013: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=83;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd210014: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=76;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd210015: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=85;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd210016: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd210017: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd210159: begin  
rid<=1;
end
19'd210160: begin  
end
19'd210161: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd210162: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd210163: begin  
rid<=0;
end
19'd210301: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=71;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5120;
 end   
19'd210302: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=36;
   mapp<=15;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4219;
 end   
19'd210303: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=19;
   mapp<=43;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7180;
 end   
19'd210304: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=84;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=9642;
 end   
19'd210305: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=57;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=7396;
 end   
19'd210306: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=84;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6915;
 end   
19'd210307: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=15;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=2702;
 end   
19'd210308: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=19;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=4650;
 end   
19'd210309: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=47;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=6618;
 end   
19'd210310: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd210311: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd210312: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=79;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=25732;
 end   
19'd210313: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=95;
   mapp<=61;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=21935;
 end   
19'd210314: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=97;
   mapp<=99;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=26472;
 end   
19'd210315: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=36;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=29489;
 end   
19'd210316: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=83;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=32389;
 end   
19'd210317: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=94;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=29665;
 end   
19'd210318: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=98;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=22251;
 end   
19'd210319: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=62;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=22327;
 end   
19'd210320: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=61;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=21284;
 end   
19'd210321: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd210322: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd210323: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd210465: begin  
rid<=1;
end
19'd210466: begin  
end
19'd210467: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd210468: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd210469: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd210470: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd210471: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd210472: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd210473: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd210474: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd210475: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd210476: begin  
rid<=0;
end
19'd210601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=54;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10363;
 end   
19'd210602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=72;
   mapp<=73;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12816;
 end   
19'd210603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=40;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd210604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=93;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd210605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=15;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd210606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=7;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd210607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd210608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=22;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=15947;
 end   
19'd210609: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=20;
   mapp<=42;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18862;
 end   
19'd210610: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=4;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd210611: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=47;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd210612: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=4;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd210613: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=1;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd210614: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd210615: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd210757: begin  
rid<=1;
end
19'd210758: begin  
end
19'd210759: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd210760: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd210761: begin  
rid<=0;
end
19'd210901: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=41;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=30961;
 end   
19'd210902: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=97;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=29129;
 end   
19'd210903: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=51;
   mapp<=98;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=31480;
 end   
19'd210904: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=61;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd210905: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=42;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd210906: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=83;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd210907: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=62;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd210908: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=88;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd210909: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=96;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd210910: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=85;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd210911: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=49;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=40755;
 end   
19'd210912: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=10;
   mapp<=51;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=38554;
 end   
19'd210913: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=23;
   mapp<=24;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=45013;
 end   
19'd210914: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=92;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd210915: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=72;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd210916: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=66;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd210917: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=8;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd210918: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=19;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd210919: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd210920: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd210921: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd211063: begin  
rid<=1;
end
19'd211064: begin  
end
19'd211065: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd211066: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd211067: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd211068: begin  
rid<=0;
end
19'd211201: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=32;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11918;
 end   
19'd211202: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=1;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd211203: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=44;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd211204: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=55;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd211205: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=54;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd211206: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=26;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=23532;
 end   
19'd211207: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=51;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd211208: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=5;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd211209: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=98;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd211210: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=56;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd211211: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd211353: begin  
rid<=1;
end
19'd211354: begin  
end
19'd211355: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd211356: begin  
rid<=0;
end
19'd211501: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=74;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12767;
 end   
19'd211502: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=13;
   mapp<=20;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12704;
 end   
19'd211503: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=44;
   mapp<=25;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=15074;
 end   
19'd211504: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=51;
   mapp<=58;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=14797;
 end   
19'd211505: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=3;
   mapp<=61;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=11502;
 end   
19'd211506: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=39;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd211507: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=56;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd211508: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=39;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd211509: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=61;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd211510: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=28;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd211511: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=10;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd211512: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=99;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=22985;
 end   
19'd211513: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=11;
   mapp<=19;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=24151;
 end   
19'd211514: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=77;
   mapp<=53;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=22635;
 end   
19'd211515: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=24;
   mapp<=13;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=26341;
 end   
19'd211516: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=19;
   mapp<=98;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=23351;
 end   
19'd211517: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=69;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd211518: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=2;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd211519: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=32;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd211520: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=54;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd211521: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=82;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd211522: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=93;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd211523: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd211665: begin  
rid<=1;
end
19'd211666: begin  
end
19'd211667: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd211668: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd211669: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd211670: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd211671: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd211672: begin  
rid<=0;
end
19'd211801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=92;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4228;
 end   
19'd211802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=14;
   mapp<=26;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1560;
 end   
19'd211803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd211804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=59;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5729;
 end   
19'd211805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=3;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=2013;
 end   
19'd211806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=8;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd211807: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd211949: begin  
rid<=1;
end
19'd211950: begin  
end
19'd211951: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd211952: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd211953: begin  
rid<=0;
end
19'd212101: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=35;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=911;
 end   
19'd212102: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=1;
   mapp<=1;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=141;
 end   
19'd212103: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=96;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3444;
 end   
19'd212104: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=64;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=2311;
 end   
19'd212105: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=41;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1516;
 end   
19'd212106: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=41;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=1584;
 end   
19'd212107: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=99;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=3532;
 end   
19'd212108: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=7;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=380;
 end   
19'd212109: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=65;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=2356;
 end   
19'd212110: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=1;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=194;
 end   
19'd212111: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd212112: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=60;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=13991;
 end   
19'd212113: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=90;
   mapp<=90;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12921;
 end   
19'd212114: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=82;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=13944;
 end   
19'd212115: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=62;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=9001;
 end   
19'd212116: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=33;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=6826;
 end   
19'd212117: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=37;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=8934;
 end   
19'd212118: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=57;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=7852;
 end   
19'd212119: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=10;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=3950;
 end   
19'd212120: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=33;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=5146;
 end   
19'd212121: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=9;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=6404;
 end   
19'd212122: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd212123: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd212265: begin  
rid<=1;
end
19'd212266: begin  
end
19'd212267: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd212268: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd212269: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd212270: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd212271: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd212272: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd212273: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd212274: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd212275: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd212276: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd212277: begin  
rid<=0;
end
19'd212401: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=70;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2030;
 end   
19'd212402: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=27;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1900;
 end   
19'd212403: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=85;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5970;
 end   
19'd212404: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=95;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6680;
 end   
19'd212405: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=45;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3190;
 end   
19'd212406: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=15;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=3350;
 end   
19'd212407: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=2425;
 end   
19'd212408: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=29;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=6405;
 end   
19'd212409: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=15;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6905;
 end   
19'd212410: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=1;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=3205;
 end   
19'd212411: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd212553: begin  
rid<=1;
end
19'd212554: begin  
end
19'd212555: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd212556: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd212557: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd212558: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd212559: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd212560: begin  
rid<=0;
end
19'd212701: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=47;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6251;
 end   
19'd212702: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=74;
   mapp<=47;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8324;
 end   
19'd212703: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=84;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd212704: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=88;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=11810;
 end   
19'd212705: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=63;
   mapp<=17;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=11979;
 end   
19'd212706: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=26;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd212707: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd212849: begin  
rid<=1;
end
19'd212850: begin  
end
19'd212851: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd212852: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd212853: begin  
rid<=0;
end
19'd213001: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=5;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=485;
 end   
19'd213002: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=52;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=270;
 end   
19'd213003: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=40;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=220;
 end   
19'd213004: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=11;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=760;
 end   
19'd213005: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=57;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=897;
 end   
19'd213006: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=49;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=759;
 end   
19'd213007: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd213149: begin  
rid<=1;
end
19'd213150: begin  
end
19'd213151: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd213152: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd213153: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd213154: begin  
rid<=0;
end
19'd213301: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=6;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=21994;
 end   
19'd213302: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=95;
   mapp<=76;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=20229;
 end   
19'd213303: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=98;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd213304: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=40;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd213305: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=8;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd213306: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=47;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd213307: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=50;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd213308: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd213309: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=59;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=36157;
 end   
19'd213310: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=60;
   mapp<=24;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=35570;
 end   
19'd213311: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=90;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd213312: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=21;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd213313: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=53;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd213314: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=21;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd213315: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=43;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd213316: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=80;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd213317: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd213459: begin  
rid<=1;
end
19'd213460: begin  
end
19'd213461: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd213462: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd213463: begin  
rid<=0;
end
19'd213601: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=89;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1780;
 end   
19'd213602: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=63;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1270;
 end   
19'd213603: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=53;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=2363;
 end   
19'd213604: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=76;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=2106;
 end   
19'd213605: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd213747: begin  
rid<=1;
end
19'd213748: begin  
end
19'd213749: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd213750: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd213751: begin  
rid<=0;
end
19'd213901: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=81;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5944;
 end   
19'd213902: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=5;
   mapp<=71;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6461;
 end   
19'd213903: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=86;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9291;
 end   
19'd213904: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=47;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=9237;
 end   
19'd213905: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=84;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=12226;
 end   
19'd213906: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=90;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=10094;
 end   
19'd213907: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=54;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=5703;
 end   
19'd213908: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=27;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd213909: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=37;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12160;
 end   
19'd213910: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=69;
   mapp<=74;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8901;
 end   
19'd213911: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=5;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=11513;
 end   
19'd213912: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=28;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=11335;
 end   
19'd213913: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=17;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=17768;
 end   
19'd213914: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=68;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=13096;
 end   
19'd213915: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=13;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=13345;
 end   
19'd213916: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=98;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd213917: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd214059: begin  
rid<=1;
end
19'd214060: begin  
end
19'd214061: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd214062: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd214063: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd214064: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd214065: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd214066: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd214067: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd214068: begin  
rid<=0;
end
19'd214201: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=90;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=17658;
 end   
19'd214202: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=76;
   mapp<=64;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15417;
 end   
19'd214203: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=55;
   mapp<=53;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=14134;
 end   
19'd214204: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=99;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd214205: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=34;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd214206: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=7;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd214207: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd214208: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd214209: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=59;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=37508;
 end   
19'd214210: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=77;
   mapp<=69;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=34056;
 end   
19'd214211: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=41;
   mapp<=12;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=33550;
 end   
19'd214212: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=83;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd214213: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=61;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd214214: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=96;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd214215: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd214216: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd214217: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd214359: begin  
rid<=1;
end
19'd214360: begin  
end
19'd214361: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd214362: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd214363: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd214364: begin  
rid<=0;
end
19'd214501: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=88;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=19406;
 end   
19'd214502: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=75;
   mapp<=62;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=17544;
 end   
19'd214503: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=78;
   mapp<=82;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=13326;
 end   
19'd214504: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=76;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7795;
 end   
19'd214505: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=5;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2481;
 end   
19'd214506: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=9;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=3755;
 end   
19'd214507: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=17;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=5783;
 end   
19'd214508: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd214509: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd214510: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=71;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=25177;
 end   
19'd214511: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=76;
   mapp<=20;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=25158;
 end   
19'd214512: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=38;
   mapp<=39;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=24151;
 end   
19'd214513: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=85;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=20328;
 end   
19'd214514: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=42;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=14279;
 end   
19'd214515: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=87;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=16734;
 end   
19'd214516: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=58;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=15259;
 end   
19'd214517: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd214518: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd214519: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd214661: begin  
rid<=1;
end
19'd214662: begin  
end
19'd214663: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd214664: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd214665: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd214666: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd214667: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd214668: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd214669: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd214670: begin  
rid<=0;
end
19'd214801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=46;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2208;
 end   
19'd214802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=14;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=654;
 end   
19'd214803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=51;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2366;
 end   
19'd214804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=36;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1686;
 end   
19'd214805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=41;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1926;
 end   
19'd214806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=50;
 end   
19'd214807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=64;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=3004;
 end   
19'd214808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=33;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5475;
 end   
19'd214809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=3195;
 end   
19'd214810: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=68;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=4610;
 end   
19'd214811: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=28;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=2610;
 end   
19'd214812: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=91;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=4929;
 end   
19'd214813: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=92;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=3086;
 end   
19'd214814: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=80;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=5644;
 end   
19'd214815: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd214957: begin  
rid<=1;
end
19'd214958: begin  
end
19'd214959: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd214960: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd214961: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd214962: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd214963: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd214964: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd214965: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd214966: begin  
rid<=0;
end
19'd215101: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=55;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4275;
 end   
19'd215102: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=20;
   mapp<=24;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2614;
 end   
19'd215103: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=51;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4379;
 end   
19'd215104: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=35;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd215105: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=99;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=9102;
 end   
19'd215106: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=32;
   mapp<=24;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=4982;
 end   
19'd215107: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=44;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=6351;
 end   
19'd215108: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=7;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd215109: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd215251: begin  
rid<=1;
end
19'd215252: begin  
end
19'd215253: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd215254: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd215255: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd215256: begin  
rid<=0;
end
19'd215401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=97;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11834;
 end   
19'd215402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=48;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10091;
 end   
19'd215403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=14;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6130;
 end   
19'd215404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=99;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=14049;
 end   
19'd215405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=92;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=11604;
 end   
19'd215406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=55;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=8841;
 end   
19'd215407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=72;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=8388;
 end   
19'd215408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd215409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=15;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=13892;
 end   
19'd215410: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=81;
   mapp<=8;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=10778;
 end   
19'd215411: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=7;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=8341;
 end   
19'd215412: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=26;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=21648;
 end   
19'd215413: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=89;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=13668;
 end   
19'd215414: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=9;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=12621;
 end   
19'd215415: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=45;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=16920;
 end   
19'd215416: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd215417: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd215559: begin  
rid<=1;
end
19'd215560: begin  
end
19'd215561: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd215562: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd215563: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd215564: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd215565: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd215566: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd215567: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd215568: begin  
rid<=0;
end
19'd215701: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=67;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=15967;
 end   
19'd215702: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=38;
   mapp<=17;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=19216;
 end   
19'd215703: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=15;
   mapp<=48;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=19502;
 end   
19'd215704: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=47;
   mapp<=14;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=16277;
 end   
19'd215705: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=73;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd215706: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=86;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd215707: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=58;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd215708: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=48;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd215709: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd215710: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd215711: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd215712: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=92;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=43348;
 end   
19'd215713: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=80;
   mapp<=36;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=46900;
 end   
19'd215714: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=17;
   mapp<=95;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=48151;
 end   
19'd215715: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=95;
   mapp<=52;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=40451;
 end   
19'd215716: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=40;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd215717: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=14;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd215718: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=29;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd215719: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=84;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd215720: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd215721: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd215722: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd215723: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd215865: begin  
rid<=1;
end
19'd215866: begin  
end
19'd215867: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd215868: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd215869: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd215870: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd215871: begin  
rid<=0;
end
19'd216001: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=4;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8229;
 end   
19'd216002: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=63;
   mapp<=53;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11330;
 end   
19'd216003: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=66;
   mapp<=67;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=13313;
 end   
19'd216004: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=5;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd216005: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=86;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd216006: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=54;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd216007: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=39;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=19152;
 end   
19'd216008: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=5;
   mapp<=94;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=30396;
 end   
19'd216009: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=81;
   mapp<=69;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=28838;
 end   
19'd216010: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=43;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd216011: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=98;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd216012: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=26;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd216013: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd216155: begin  
rid<=1;
end
19'd216156: begin  
end
19'd216157: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd216158: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd216159: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd216160: begin  
rid<=0;
end
19'd216301: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=95;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13984;
 end   
19'd216302: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=6;
   mapp<=69;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11055;
 end   
19'd216303: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=47;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9621;
 end   
19'd216304: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=60;
   mapp<=70;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=12042;
 end   
19'd216305: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd216306: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd216307: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd216308: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=33;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=31856;
 end   
19'd216309: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=95;
   mapp<=81;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=28461;
 end   
19'd216310: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=28;
   mapp<=94;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=26138;
 end   
19'd216311: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=49;
   mapp<=90;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=24898;
 end   
19'd216312: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd216313: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd216314: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd216315: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd216457: begin  
rid<=1;
end
19'd216458: begin  
end
19'd216459: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd216460: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd216461: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd216462: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd216463: begin  
rid<=0;
end
19'd216601: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=74;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14537;
 end   
19'd216602: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=83;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10110;
 end   
19'd216603: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=16;
   mapp<=51;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9541;
 end   
19'd216604: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=83;
   mapp<=56;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6194;
 end   
19'd216605: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=38;
   mapp<=1;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5371;
 end   
19'd216606: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=4;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7485;
 end   
19'd216607: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=6;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=13172;
 end   
19'd216608: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=63;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd216609: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=63;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd216610: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=80;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd216611: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd216612: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=6;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=21872;
 end   
19'd216613: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=71;
   mapp<=34;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=16190;
 end   
19'd216614: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=3;
   mapp<=56;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=18541;
 end   
19'd216615: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=64;
   mapp<=73;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=18800;
 end   
19'd216616: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=1;
   mapp<=75;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=18263;
 end   
19'd216617: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=30;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=23289;
 end   
19'd216618: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=61;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=25948;
 end   
19'd216619: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=85;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd216620: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=30;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd216621: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=90;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd216622: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=21;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd216623: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd216765: begin  
rid<=1;
end
19'd216766: begin  
end
19'd216767: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd216768: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd216769: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd216770: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd216771: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd216772: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd216773: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd216774: begin  
rid<=0;
end
19'd216901: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=26;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12410;
 end   
19'd216902: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=27;
   mapp<=44;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12176;
 end   
19'd216903: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=80;
   mapp<=39;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11819;
 end   
19'd216904: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=79;
   mapp<=94;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=15076;
 end   
19'd216905: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=31;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=11977;
 end   
19'd216906: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=73;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=9859;
 end   
19'd216907: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=75;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=11103;
 end   
19'd216908: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd216909: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd216910: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd216911: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=57;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=24435;
 end   
19'd216912: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=67;
   mapp<=92;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=23870;
 end   
19'd216913: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=23;
   mapp<=64;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=23674;
 end   
19'd216914: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=94;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=27168;
 end   
19'd216915: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=83;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=21873;
 end   
19'd216916: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=51;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=20043;
 end   
19'd216917: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=76;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=23134;
 end   
19'd216918: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd216919: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd216920: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd216921: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd217063: begin  
rid<=1;
end
19'd217064: begin  
end
19'd217065: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd217066: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd217067: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd217068: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd217069: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd217070: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd217071: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd217072: begin  
rid<=0;
end
19'd217201: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=52;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16275;
 end   
19'd217202: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=6;
   mapp<=65;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=18988;
 end   
19'd217203: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=50;
   mapp<=77;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=22250;
 end   
19'd217204: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=62;
   mapp<=51;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=21214;
 end   
19'd217205: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=77;
   mapp<=43;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=18238;
 end   
19'd217206: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=82;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd217207: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=73;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd217208: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd217209: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=20;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd217210: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=1;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd217211: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=35;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=27377;
 end   
19'd217212: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=19;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=31589;
 end   
19'd217213: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=16;
   mapp<=80;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=37474;
 end   
19'd217214: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=40;
   mapp<=66;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=38289;
 end   
19'd217215: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=42;
   mapp<=37;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=33886;
 end   
19'd217216: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=91;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd217217: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd217218: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd217219: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=35;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd217220: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=14;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd217221: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd217363: begin  
rid<=1;
end
19'd217364: begin  
end
19'd217365: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd217366: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd217367: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd217368: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd217369: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd217370: begin  
rid<=0;
end
19'd217501: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=67;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12637;
 end   
19'd217502: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=45;
   mapp<=18;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15115;
 end   
19'd217503: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=13;
   mapp<=18;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8126;
 end   
19'd217504: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=57;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd217505: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=19;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd217506: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=76;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd217507: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=8;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd217508: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=48;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd217509: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd217510: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=97;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd217511: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=73;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=31099;
 end   
19'd217512: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=94;
   mapp<=10;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=31687;
 end   
19'd217513: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=29;
   mapp<=71;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=27518;
 end   
19'd217514: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=33;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd217515: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=75;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd217516: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=62;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd217517: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=88;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd217518: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=15;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd217519: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd217520: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=30;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd217521: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd217663: begin  
rid<=1;
end
19'd217664: begin  
end
19'd217665: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd217666: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd217667: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd217668: begin  
rid<=0;
end
19'd217801: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=10;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=375;
 end   
19'd217802: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=9;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=483;
 end   
19'd217803: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=47;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=940;
 end   
19'd217804: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=50;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=728;
 end   
19'd217805: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=22;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=719;
 end   
19'd217806: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=51;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=821;
 end   
19'd217807: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=29;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=827;
 end   
19'd217808: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=53;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=1023;
 end   
19'd217809: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd217810: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=74;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7153;
 end   
19'd217811: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=1;
   mapp<=44;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=3812;
 end   
19'd217812: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=73;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=6379;
 end   
19'd217813: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=37;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=3493;
 end   
19'd217814: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=27;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=2793;
 end   
19'd217815: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=76;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=6514;
 end   
19'd217816: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=69;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=6017;
 end   
19'd217817: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=84;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=7273;
 end   
19'd217818: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd217819: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd217961: begin  
rid<=1;
end
19'd217962: begin  
end
19'd217963: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd217964: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd217965: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd217966: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd217967: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd217968: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd217969: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd217970: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd217971: begin  
rid<=0;
end
19'd218101: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=5;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=85;
 end   
19'd218102: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=16;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=90;
 end   
19'd218103: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=84;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=440;
 end   
19'd218104: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=84;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=450;
 end   
19'd218105: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=41;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=1561;
 end   
19'd218106: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=59;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=2509;
 end   
19'd218107: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=9;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=809;
 end   
19'd218108: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=27;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=1557;
 end   
19'd218109: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd218251: begin  
rid<=1;
end
19'd218252: begin  
end
19'd218253: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd218254: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd218255: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd218256: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd218257: begin  
rid<=0;
end
19'd218401: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=43;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=28650;
 end   
19'd218402: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=71;
   mapp<=66;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=36722;
 end   
19'd218403: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=86;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd218404: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=80;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd218405: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=85;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd218406: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=5;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd218407: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=67;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd218408: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=34;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd218409: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=54;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd218410: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd218411: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=65;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=50187;
 end   
19'd218412: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=10;
   mapp<=57;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=57706;
 end   
19'd218413: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=22;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd218414: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=43;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd218415: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=74;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd218416: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=8;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd218417: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=42;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd218418: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=29;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd218419: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=82;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd218420: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd218421: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd218563: begin  
rid<=1;
end
19'd218564: begin  
end
19'd218565: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd218566: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd218567: begin  
rid<=0;
end
19'd218701: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=52;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13303;
 end   
19'd218702: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=32;
   mapp<=62;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15714;
 end   
19'd218703: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=97;
   mapp<=99;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12508;
 end   
19'd218704: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd218705: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd218706: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=72;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=21143;
 end   
19'd218707: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=77;
   mapp<=12;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=25152;
 end   
19'd218708: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=50;
   mapp<=62;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=27574;
 end   
19'd218709: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd218710: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd218711: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd218853: begin  
rid<=1;
end
19'd218854: begin  
end
19'd218855: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd218856: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd218857: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd218858: begin  
rid<=0;
end
19'd219001: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=26;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13832;
 end   
19'd219002: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=8;
   mapp<=64;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=18084;
 end   
19'd219003: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=35;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd219004: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=42;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd219005: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=67;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd219006: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=54;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd219007: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=47;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd219008: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=5;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd219009: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=84;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd219010: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=53;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd219011: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=46;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=37171;
 end   
19'd219012: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=20;
   mapp<=41;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=38309;
 end   
19'd219013: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=97;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd219014: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=71;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd219015: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=46;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd219016: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=81;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd219017: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=11;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd219018: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=28;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd219019: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=46;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd219020: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=90;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd219021: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd219163: begin  
rid<=1;
end
19'd219164: begin  
end
19'd219165: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd219166: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd219167: begin  
rid<=0;
end
19'd219301: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=72;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14453;
 end   
19'd219302: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=38;
   mapp<=88;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=19757;
 end   
19'd219303: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=70;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd219304: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=76;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd219305: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=5;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd219306: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=32;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd219307: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=29;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd219308: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=19;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd219309: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd219310: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=61;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=47190;
 end   
19'd219311: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=43;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=57044;
 end   
19'd219312: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=69;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd219313: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=4;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd219314: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=84;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd219315: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=97;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd219316: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=71;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd219317: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=84;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd219318: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd219319: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd219461: begin  
rid<=1;
end
19'd219462: begin  
end
19'd219463: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd219464: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd219465: begin  
rid<=0;
end
19'd219601: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=54;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1404;
 end   
19'd219602: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=87;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4708;
 end   
19'd219603: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=48;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2612;
 end   
19'd219604: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=31;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=4101;
 end   
19'd219605: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=9;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=4987;
 end   
19'd219606: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=7;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=2829;
 end   
19'd219607: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd219749: begin  
rid<=1;
end
19'd219750: begin  
end
19'd219751: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd219752: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd219753: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd219754: begin  
rid<=0;
end
19'd219901: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=88;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9197;
 end   
19'd219902: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=67;
   mapp<=60;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9146;
 end   
19'd219903: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=29;
   mapp<=45;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7054;
 end   
19'd219904: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=29;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5456;
 end   
19'd219905: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=39;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4684;
 end   
19'd219906: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=9;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=4221;
 end   
19'd219907: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=21;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=8436;
 end   
19'd219908: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=68;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=11944;
 end   
19'd219909: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=68;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=9610;
 end   
19'd219910: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd219911: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd219912: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=78;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16326;
 end   
19'd219913: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=41;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18278;
 end   
19'd219914: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=58;
   mapp<=50;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15572;
 end   
19'd219915: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=32;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=15451;
 end   
19'd219916: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=57;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=14751;
 end   
19'd219917: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=89;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=15979;
 end   
19'd219918: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=34;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=18901;
 end   
19'd219919: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=59;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=24013;
 end   
19'd219920: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=93;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=19795;
 end   
19'd219921: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd219922: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd219923: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd220065: begin  
rid<=1;
end
19'd220066: begin  
end
19'd220067: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd220068: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd220069: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd220070: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd220071: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd220072: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd220073: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd220074: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd220075: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd220076: begin  
rid<=0;
end
19'd220201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=17;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3726;
 end   
19'd220202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=13;
   mapp<=29;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2511;
 end   
19'd220203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=51;
   mapp<=57;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2093;
 end   
19'd220204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=12;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=2540;
 end   
19'd220205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=7;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2092;
 end   
19'd220206: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=35;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6069;
 end   
19'd220207: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=15;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=4310;
 end   
19'd220208: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=82;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=5977;
 end   
19'd220209: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=26;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd220210: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=53;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd220211: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=87;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12400;
 end   
19'd220212: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=31;
   mapp<=52;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8445;
 end   
19'd220213: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=48;
   mapp<=13;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=11248;
 end   
19'd220214: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=88;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=14369;
 end   
19'd220215: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=79;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=14035;
 end   
19'd220216: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=93;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=19282;
 end   
19'd220217: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=97;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=17520;
 end   
19'd220218: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=99;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=17021;
 end   
19'd220219: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=68;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd220220: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=14;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd220221: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd220363: begin  
rid<=1;
end
19'd220364: begin  
end
19'd220365: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd220366: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd220367: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd220368: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd220369: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd220370: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd220371: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd220372: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd220373: begin  
rid<=0;
end
19'd220501: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=38;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5983;
 end   
19'd220502: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=87;
   mapp<=34;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7709;
 end   
19'd220503: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=71;
   mapp<=41;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11306;
 end   
19'd220504: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd220505: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd220506: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=73;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14093;
 end   
19'd220507: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=66;
   mapp<=82;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=15975;
 end   
19'd220508: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=12;
   mapp<=18;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=18734;
 end   
19'd220509: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd220510: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd220511: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd220653: begin  
rid<=1;
end
19'd220654: begin  
end
19'd220655: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd220656: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd220657: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd220658: begin  
rid<=0;
end
19'd220801: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=5;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1159;
 end   
19'd220802: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=49;
   mapp<=21;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3741;
 end   
19'd220803: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=74;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2742;
 end   
19'd220804: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=48;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=2818;
 end   
19'd220805: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=52;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4318;
 end   
19'd220806: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=82;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=4135;
 end   
19'd220807: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=75;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=3718;
 end   
19'd220808: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=67;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=5207;
 end   
19'd220809: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=98;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=2824;
 end   
19'd220810: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=46;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=4975;
 end   
19'd220811: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd220812: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=15;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=1789;
 end   
19'd220813: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=25;
   mapp<=15;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=5641;
 end   
19'd220814: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=67;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=5972;
 end   
19'd220815: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=89;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6153;
 end   
19'd220816: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=80;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=7343;
 end   
19'd220817: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=73;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=6755;
 end   
19'd220818: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=61;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=6883;
 end   
19'd220819: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=90;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=7032;
 end   
19'd220820: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=19;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=3334;
 end   
19'd220821: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=9;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=6910;
 end   
19'd220822: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd220823: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd220965: begin  
rid<=1;
end
19'd220966: begin  
end
19'd220967: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd220968: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd220969: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd220970: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd220971: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd220972: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd220973: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd220974: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd220975: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd220976: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd220977: begin  
rid<=0;
end
19'd221101: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=57;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3078;
 end   
19'd221102: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5425;
 end   
19'd221103: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=7;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=419;
 end   
19'd221104: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=37;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=2139;
 end   
19'd221105: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=83;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4771;
 end   
19'd221106: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=99;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=9315;
 end   
19'd221107: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=5623;
 end   
19'd221108: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=96;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=9923;
 end   
19'd221109: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=90;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=11049;
 end   
19'd221110: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=16;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=6355;
 end   
19'd221111: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd221253: begin  
rid<=1;
end
19'd221254: begin  
end
19'd221255: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd221256: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd221257: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd221258: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd221259: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd221260: begin  
rid<=0;
end
19'd221401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=45;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6999;
 end   
19'd221402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=84;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4925;
 end   
19'd221403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=4;
   mapp<=39;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5268;
 end   
19'd221404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=61;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5982;
 end   
19'd221405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=27;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=7397;
 end   
19'd221406: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=64;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd221407: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=60;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd221408: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=80;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16311;
 end   
19'd221409: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=6;
   mapp<=12;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8077;
 end   
19'd221410: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=51;
   mapp<=40;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=13578;
 end   
19'd221411: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=50;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=13338;
 end   
19'd221412: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=78;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=15793;
 end   
19'd221413: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=48;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd221414: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=20;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd221415: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd221557: begin  
rid<=1;
end
19'd221558: begin  
end
19'd221559: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd221560: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd221561: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd221562: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd221563: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd221564: begin  
rid<=0;
end
19'd221701: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=35;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1400;
 end   
19'd221702: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=42;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1690;
 end   
19'd221703: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=9;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=380;
 end   
19'd221704: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=43;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=2475;
 end   
19'd221705: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=95;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=4065;
 end   
19'd221706: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=57;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=1805;
 end   
19'd221707: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd221849: begin  
rid<=1;
end
19'd221850: begin  
end
19'd221851: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd221852: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd221853: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd221854: begin  
rid<=0;
end
19'd222001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=31;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4221;
 end   
19'd222002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=18;
   mapp<=91;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4883;
 end   
19'd222003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=18;
   mapp<=35;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2653;
 end   
19'd222004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=79;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3829;
 end   
19'd222005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=7;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2651;
 end   
19'd222006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=68;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=3616;
 end   
19'd222007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=65;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=4037;
 end   
19'd222008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=16;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=3554;
 end   
19'd222009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=93;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=5699;
 end   
19'd222010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd222011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd222012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=85;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=18382;
 end   
19'd222013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=83;
   mapp<=78;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=14042;
 end   
19'd222014: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=29;
   mapp<=13;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=8633;
 end   
19'd222015: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=50;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=10908;
 end   
19'd222016: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=25;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=9196;
 end   
19'd222017: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=26;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=14417;
 end   
19'd222018: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=78;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=16755;
 end   
19'd222019: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=73;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=9958;
 end   
19'd222020: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=1;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=8523;
 end   
19'd222021: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd222022: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd222023: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd222165: begin  
rid<=1;
end
19'd222166: begin  
end
19'd222167: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd222168: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd222169: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd222170: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd222171: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd222172: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd222173: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd222174: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd222175: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd222176: begin  
rid<=0;
end
19'd222301: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=68;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4556;
 end   
19'd222302: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=47;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3159;
 end   
19'd222303: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=43;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2901;
 end   
19'd222304: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=47;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3179;
 end   
19'd222305: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=57;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3859;
 end   
19'd222306: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=11;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=787;
 end   
19'd222307: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=73;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=4951;
 end   
19'd222308: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=97;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=6569;
 end   
19'd222309: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=49;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=3363;
 end   
19'd222310: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=37;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=2569;
 end   
19'd222311: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=95;
   mapp<=0;
   pp<=100;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[10]<=6465;
 end   
19'd222312: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=7;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=4696;
 end   
19'd222313: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=68;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=4519;
 end   
19'd222314: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=47;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=3841;
 end   
19'd222315: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=3179;
 end   
19'd222316: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=61;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=5079;
 end   
19'd222317: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=33;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=1447;
 end   
19'd222318: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=16;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=5271;
 end   
19'd222319: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=93;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=8429;
 end   
19'd222320: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=7;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=3503;
 end   
19'd222321: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=50;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=3569;
 end   
19'd222322: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=75;
   mapp<=0;
   pp<=100;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[10]<=7965;
 end   
19'd222323: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd222465: begin  
rid<=1;
end
19'd222466: begin  
end
19'd222467: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd222468: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd222469: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd222470: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd222471: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd222472: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd222473: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd222474: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd222475: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd222476: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd222477: begin  
check0<=expctdoutput[10]-outcheck0;
end
19'd222478: begin  
rid<=0;
end
19'd222601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=14;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=18333;
 end   
19'd222602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=85;
   mapp<=78;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=14989;
 end   
19'd222603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=31;
   mapp<=86;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7022;
 end   
19'd222604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=52;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd222605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=10;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd222606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=5;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd222607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=74;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd222608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd222609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd222610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=33;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=33699;
 end   
19'd222611: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=57;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=30808;
 end   
19'd222612: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=47;
   mapp<=50;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=23392;
 end   
19'd222613: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=51;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd222614: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=93;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd222615: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=34;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd222616: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=61;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd222617: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd222618: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd222619: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd222761: begin  
rid<=1;
end
19'd222762: begin  
end
19'd222763: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd222764: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd222765: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd222766: begin  
rid<=0;
end
19'd222901: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=63;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=21084;
 end   
19'd222902: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=66;
   mapp<=79;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=22957;
 end   
19'd222903: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=84;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd222904: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=47;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd222905: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=87;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd222906: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=56;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd222907: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd222908: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=49;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=40329;
 end   
19'd222909: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=41;
   mapp<=55;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=41026;
 end   
19'd222910: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=33;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd222911: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=29;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd222912: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=61;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd222913: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=92;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd222914: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd222915: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd223057: begin  
rid<=1;
end
19'd223058: begin  
end
19'd223059: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd223060: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd223061: begin  
rid<=0;
end
19'd223201: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=90;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16740;
 end   
19'd223202: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=84;
   mapp<=57;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=13284;
 end   
19'd223203: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=34;
   mapp<=81;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=14694;
 end   
19'd223204: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=58;
   mapp<=36;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=8854;
 end   
19'd223205: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd223206: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd223207: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd223208: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=74;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=28295;
 end   
19'd223209: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=86;
   mapp<=6;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=27732;
 end   
19'd223210: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=17;
   mapp<=53;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=27167;
 end   
19'd223211: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=89;
   mapp<=74;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=24052;
 end   
19'd223212: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd223213: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd223214: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd223215: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd223357: begin  
rid<=1;
end
19'd223358: begin  
end
19'd223359: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd223360: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd223361: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd223362: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd223363: begin  
rid<=0;
end
19'd223501: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=89;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6853;
 end   
19'd223502: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=47;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4193;
 end   
19'd223503: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=1;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=109;
 end   
19'd223504: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=61;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5459;
 end   
19'd223505: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=29;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2621;
 end   
19'd223506: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=3;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=317;
 end   
19'd223507: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=92;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=8248;
 end   
19'd223508: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=25;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=2295;
 end   
19'd223509: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=99;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=8891;
 end   
19'd223510: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=92;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12741;
 end   
19'd223511: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=88;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12289;
 end   
19'd223512: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=95;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=8849;
 end   
19'd223513: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=67;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=11623;
 end   
19'd223514: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=22;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=4645;
 end   
19'd223515: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=70;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=6757;
 end   
19'd223516: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=73;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=14964;
 end   
19'd223517: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=2;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=2479;
 end   
19'd223518: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=63;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=14687;
 end   
19'd223519: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd223661: begin  
rid<=1;
end
19'd223662: begin  
end
19'd223663: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd223664: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd223665: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd223666: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd223667: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd223668: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd223669: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd223670: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd223671: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd223672: begin  
rid<=0;
end
19'd223801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=88;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16914;
 end   
19'd223802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=46;
   mapp<=34;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15828;
 end   
19'd223803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=56;
   mapp<=99;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=18510;
 end   
19'd223804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=54;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd223805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=60;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd223806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=6;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd223807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=51;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd223808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=28;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd223809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=74;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd223810: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=97;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=43682;
 end   
19'd223811: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=70;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=44463;
 end   
19'd223812: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=89;
   mapp<=63;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=37140;
 end   
19'd223813: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=60;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd223814: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=93;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd223815: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=73;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd223816: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=19;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd223817: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=54;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd223818: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=10;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd223819: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd223961: begin  
rid<=1;
end
19'd223962: begin  
end
19'd223963: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd223964: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd223965: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd223966: begin  
rid<=0;
end
19'd224101: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=75;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11821;
 end   
19'd224102: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=44;
   mapp<=98;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=13849;
 end   
19'd224103: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=56;
   mapp<=66;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11435;
 end   
19'd224104: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=38;
   mapp<=51;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=12077;
 end   
19'd224105: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=93;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=9508;
 end   
19'd224106: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=3;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=11979;
 end   
19'd224107: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=35;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=17292;
 end   
19'd224108: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd224109: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=50;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd224110: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=85;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd224111: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=84;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=27347;
 end   
19'd224112: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=64;
   mapp<=81;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=25064;
 end   
19'd224113: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=52;
   mapp<=91;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=20134;
 end   
19'd224114: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=33;
   mapp<=30;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=21485;
 end   
19'd224115: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=16;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=19302;
 end   
19'd224116: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=57;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=23902;
 end   
19'd224117: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=37;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=32317;
 end   
19'd224118: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=31;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd224119: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=99;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd224120: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=49;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd224121: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd224263: begin  
rid<=1;
end
19'd224264: begin  
end
19'd224265: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd224266: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd224267: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd224268: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd224269: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd224270: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd224271: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd224272: begin  
rid<=0;
end
19'd224401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=58;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14194;
 end   
19'd224402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=95;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=14251;
 end   
19'd224403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=94;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd224404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=73;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd224405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=56;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd224406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=62;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd224407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=23;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd224408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd224409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=63;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=37184;
 end   
19'd224410: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=86;
   mapp<=63;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=35538;
 end   
19'd224411: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=72;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd224412: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=44;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd224413: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=19;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd224414: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=66;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd224415: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=70;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd224416: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd224417: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd224559: begin  
rid<=1;
end
19'd224560: begin  
end
19'd224561: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd224562: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd224563: begin  
rid<=0;
end
19'd224701: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=24;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7830;
 end   
19'd224702: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=5;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8442;
 end   
19'd224703: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=93;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd224704: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=34;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd224705: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd224706: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=79;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=15426;
 end   
19'd224707: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=74;
   mapp<=41;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=13199;
 end   
19'd224708: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=7;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd224709: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=26;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd224710: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=0;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd224711: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd224853: begin  
rid<=1;
end
19'd224854: begin  
end
19'd224855: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd224856: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd224857: begin  
rid<=0;
end
19'd225001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=41;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9228;
 end   
19'd225002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=9;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12184;
 end   
19'd225003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=61;
   mapp<=16;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=15809;
 end   
19'd225004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=72;
   mapp<=70;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=8474;
 end   
19'd225005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=35;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd225006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=87;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd225007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=3;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd225008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd225009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=36;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16612;
 end   
19'd225010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=50;
   mapp<=21;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=26491;
 end   
19'd225011: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=2;
   mapp<=73;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=21696;
 end   
19'd225012: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=58;
   mapp<=13;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=25976;
 end   
19'd225013: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=37;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd225014: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=80;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd225015: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=11;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd225016: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd225017: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd225159: begin  
rid<=1;
end
19'd225160: begin  
end
19'd225161: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd225162: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd225163: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd225164: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd225165: begin  
rid<=0;
end
19'd225301: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=23;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=15281;
 end   
19'd225302: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=84;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=19495;
 end   
19'd225303: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=91;
   mapp<=1;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=16165;
 end   
19'd225304: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=11;
   mapp<=5;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=14841;
 end   
19'd225305: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=74;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd225306: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=36;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd225307: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=94;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd225308: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=72;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd225309: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd225310: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=45;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd225311: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=70;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=31713;
 end   
19'd225312: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=17;
   mapp<=59;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=37674;
 end   
19'd225313: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=8;
   mapp<=27;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=27837;
 end   
19'd225314: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=49;
   mapp<=69;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=32423;
 end   
19'd225315: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=70;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd225316: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=14;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd225317: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=86;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd225318: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=92;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd225319: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=1;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd225320: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=35;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd225321: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd225463: begin  
rid<=1;
end
19'd225464: begin  
end
19'd225465: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd225466: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd225467: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd225468: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd225469: begin  
rid<=0;
end
19'd225601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=82;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7585;
 end   
19'd225602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=79;
   mapp<=41;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5584;
 end   
19'd225603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=28;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9031;
 end   
19'd225604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=85;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=14584;
 end   
19'd225605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=96;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=15496;
 end   
19'd225606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=96;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=12346;
 end   
19'd225607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd225608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=24;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12065;
 end   
19'd225609: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=58;
   mapp<=64;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12166;
 end   
19'd225610: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=87;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=16107;
 end   
19'd225611: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=86;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=17228;
 end   
19'd225612: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=10;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=15794;
 end   
19'd225613: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=1;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=13124;
 end   
19'd225614: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd225615: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd225757: begin  
rid<=1;
end
19'd225758: begin  
end
19'd225759: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd225760: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd225761: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd225762: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd225763: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd225764: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd225765: begin  
rid<=0;
end
19'd225901: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=32;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1582;
 end   
19'd225902: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=5;
   mapp<=86;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=878;
 end   
19'd225903: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=8;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4350;
 end   
19'd225904: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=47;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6022;
 end   
19'd225905: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=50;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=9838;
 end   
19'd225906: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=93;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd225907: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=83;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7637;
 end   
19'd225908: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=20;
   mapp<=33;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=3102;
 end   
19'd225909: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=28;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=7259;
 end   
19'd225910: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=33;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=10246;
 end   
19'd225911: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=63;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=16474;
 end   
19'd225912: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=77;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd225913: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd226055: begin  
rid<=1;
end
19'd226056: begin  
end
19'd226057: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd226058: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd226059: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd226060: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd226061: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd226062: begin  
rid<=0;
end
19'd226201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=70;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10066;
 end   
19'd226202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=85;
   mapp<=80;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6679;
 end   
19'd226203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=32;
   mapp<=39;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3531;
 end   
19'd226204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=3;
   mapp<=66;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3945;
 end   
19'd226205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=27;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=7879;
 end   
19'd226206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=21;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7267;
 end   
19'd226207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=13;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=11033;
 end   
19'd226208: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=75;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd226209: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=41;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd226210: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=46;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd226211: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=19;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=22634;
 end   
19'd226212: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=2;
   mapp<=64;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=19497;
 end   
19'd226213: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=57;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=18867;
 end   
19'd226214: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=89;
   mapp<=80;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=18895;
 end   
19'd226215: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=35;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=17069;
 end   
19'd226216: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=40;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=16171;
 end   
19'd226217: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=46;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=22331;
 end   
19'd226218: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd226219: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=29;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd226220: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=66;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd226221: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd226363: begin  
rid<=1;
end
19'd226364: begin  
end
19'd226365: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd226366: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd226367: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd226368: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd226369: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd226370: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd226371: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd226372: begin  
rid<=0;
end
19'd226501: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=52;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=728;
 end   
19'd226502: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=98;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1382;
 end   
19'd226503: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=37;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=538;
 end   
19'd226504: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=95;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1360;
 end   
19'd226505: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=10;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=180;
 end   
19'd226506: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=7;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=148;
 end   
19'd226507: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=18;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=312;
 end   
19'd226508: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=80;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=1190;
 end   
19'd226509: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=73;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=1102;
 end   
19'd226510: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=72;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=3392;
 end   
19'd226511: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=84;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=4490;
 end   
19'd226512: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=34;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=1796;
 end   
19'd226513: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=84;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=4468;
 end   
19'd226514: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=93;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=3621;
 end   
19'd226515: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=63;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=2479;
 end   
19'd226516: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=33;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=1533;
 end   
19'd226517: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=42;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=2744;
 end   
19'd226518: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=49;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=2915;
 end   
19'd226519: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd226661: begin  
rid<=1;
end
19'd226662: begin  
end
19'd226663: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd226664: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd226665: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd226666: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd226667: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd226668: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd226669: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd226670: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd226671: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd226672: begin  
rid<=0;
end
19'd226801: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=41;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10510;
 end   
19'd226802: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=72;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7947;
 end   
19'd226803: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=55;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7963;
 end   
19'd226804: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=79;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3845;
 end   
19'd226805: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=8;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=440;
 end   
19'd226806: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=1;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=5563;
 end   
19'd226807: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=76;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=6056;
 end   
19'd226808: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=40;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=6534;
 end   
19'd226809: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd226810: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=14;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12987;
 end   
19'd226811: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=37;
   mapp<=31;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=10749;
 end   
19'd226812: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=64;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=11634;
 end   
19'd226813: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=75;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=7781;
 end   
19'd226814: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=78;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=4751;
 end   
19'd226815: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=87;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=9075;
 end   
19'd226816: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=62;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=7849;
 end   
19'd226817: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=25;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=10547;
 end   
19'd226818: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd226819: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd226961: begin  
rid<=1;
end
19'd226962: begin  
end
19'd226963: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd226964: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd226965: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd226966: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd226967: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd226968: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd226969: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd226970: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd226971: begin  
rid<=0;
end
19'd227101: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=91;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=24065;
 end   
19'd227102: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=88;
   mapp<=58;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=20173;
 end   
19'd227103: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=31;
   mapp<=68;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=21210;
 end   
19'd227104: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=85;
   mapp<=88;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=19690;
 end   
19'd227105: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=15;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd227106: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=3;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd227107: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=66;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd227108: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=23;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd227109: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=80;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd227110: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=5;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd227111: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd227112: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=76;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=37450;
 end   
19'd227113: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=67;
   mapp<=39;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=32555;
 end   
19'd227114: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=53;
   mapp<=14;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=33611;
 end   
19'd227115: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=10;
   mapp<=48;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=34839;
 end   
19'd227116: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=78;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd227117: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=1;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd227118: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=12;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd227119: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=36;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd227120: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=73;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd227121: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=19;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd227122: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=99;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd227123: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd227265: begin  
rid<=1;
end
19'd227266: begin  
end
19'd227267: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd227268: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd227269: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd227270: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd227271: begin  
rid<=0;
end
19'd227401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=80;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9580;
 end   
19'd227402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=65;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd227403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=49;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd227404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=15;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12174;
 end   
19'd227405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=9;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd227406: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=67;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd227407: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd227549: begin  
rid<=1;
end
19'd227550: begin  
end
19'd227551: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd227552: begin  
rid<=0;
end
19'd227701: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=88;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10754;
 end   
19'd227702: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=71;
   mapp<=6;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8026;
 end   
19'd227703: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=48;
   mapp<=96;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=13206;
 end   
19'd227704: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=14;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=9200;
 end   
19'd227705: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd227706: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd227707: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=32;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17070;
 end   
19'd227708: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=22;
   mapp<=26;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=10453;
 end   
19'd227709: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=77;
   mapp<=48;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=21364;
 end   
19'd227710: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=7;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=15584;
 end   
19'd227711: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd227712: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd227713: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd227855: begin  
rid<=1;
end
19'd227856: begin  
end
19'd227857: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd227858: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd227859: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd227860: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd227861: begin  
rid<=0;
end
19'd228001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=84;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12639;
 end   
19'd228002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=53;
   mapp<=99;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10605;
 end   
19'd228003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=43;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7448;
 end   
19'd228004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=72;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=8887;
 end   
19'd228005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd228006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=50;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14883;
 end   
19'd228007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=22;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=14807;
 end   
19'd228008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=16;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=8930;
 end   
19'd228009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=31;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=12417;
 end   
19'd228010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd228011: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd228153: begin  
rid<=1;
end
19'd228154: begin  
end
19'd228155: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd228156: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd228157: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd228158: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd228159: begin  
rid<=0;
end
19'd228301: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=85;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11745;
 end   
19'd228302: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=89;
   mapp<=80;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9069;
 end   
19'd228303: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=30;
   mapp<=21;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5032;
 end   
19'd228304: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=13;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=9976;
 end   
19'd228305: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=69;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=14305;
 end   
19'd228306: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd228307: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd228308: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=26;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17693;
 end   
19'd228309: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=56;
   mapp<=59;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=16007;
 end   
19'd228310: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=15;
   mapp<=74;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=11795;
 end   
19'd228311: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=84;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=13969;
 end   
19'd228312: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=9;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=19786;
 end   
19'd228313: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd228314: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd228315: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd228457: begin  
rid<=1;
end
19'd228458: begin  
end
19'd228459: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd228460: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd228461: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd228462: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd228463: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd228464: begin  
rid<=0;
end
19'd228601: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=52;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2132;
 end   
19'd228602: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=60;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2470;
 end   
19'd228603: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=15;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=635;
 end   
19'd228604: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=76;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3146;
 end   
19'd228605: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=56;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2336;
 end   
19'd228606: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=43;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=1813;
 end   
19'd228607: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=42;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=1782;
 end   
19'd228608: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=40;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=4172;
 end   
19'd228609: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=66;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=5836;
 end   
19'd228610: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=6;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=941;
 end   
19'd228611: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=98;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=8144;
 end   
19'd228612: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=71;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=5957;
 end   
19'd228613: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=40;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=3853;
 end   
19'd228614: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=70;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=5352;
 end   
19'd228615: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd228757: begin  
rid<=1;
end
19'd228758: begin  
end
19'd228759: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd228760: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd228761: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd228762: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd228763: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd228764: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd228765: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd228766: begin  
rid<=0;
end
19'd228901: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=30;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10947;
 end   
19'd228902: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=27;
   mapp<=1;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11770;
 end   
19'd228903: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=61;
   mapp<=44;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=16794;
 end   
19'd228904: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=34;
   mapp<=25;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=14929;
 end   
19'd228905: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=74;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd228906: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=95;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd228907: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=23;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd228908: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd228909: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd228910: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd228911: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=54;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=29439;
 end   
19'd228912: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=45;
   mapp<=79;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=34618;
 end   
19'd228913: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=51;
   mapp<=88;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=36488;
 end   
19'd228914: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=8;
   mapp<=93;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=32716;
 end   
19'd228915: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=85;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd228916: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=48;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd228917: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=6;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd228918: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd228919: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd228920: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd228921: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd229063: begin  
rid<=1;
end
19'd229064: begin  
end
19'd229065: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd229066: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd229067: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd229068: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd229069: begin  
rid<=0;
end
19'd229201: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=20;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1968;
 end   
19'd229202: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=7;
   mapp<=64;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1507;
 end   
19'd229203: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=31;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=850;
 end   
19'd229204: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=30;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=924;
 end   
19'd229205: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd229206: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=56;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=6322;
 end   
19'd229207: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=7;
   mapp<=86;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=6841;
 end   
19'd229208: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=74;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=5631;
 end   
19'd229209: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=91;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6601;
 end   
19'd229210: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd229211: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd229353: begin  
rid<=1;
end
19'd229354: begin  
end
19'd229355: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd229356: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd229357: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd229358: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd229359: begin  
rid<=0;
end
19'd229501: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=42;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5194;
 end   
19'd229502: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=34;
   mapp<=63;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4772;
 end   
19'd229503: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=14;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd229504: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd229505: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=35;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8389;
 end   
19'd229506: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=40;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=9360;
 end   
19'd229507: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=1;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd229508: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd229509: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd229651: begin  
rid<=1;
end
19'd229652: begin  
end
19'd229653: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd229654: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd229655: begin  
rid<=0;
end
19'd229801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=89;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16588;
 end   
19'd229802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=64;
   mapp<=84;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=16425;
 end   
19'd229803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=10;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd229804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=8;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd229805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=2;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd229806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=85;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd229807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=81;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd229808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=58;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=25984;
 end   
19'd229809: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=52;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=27569;
 end   
19'd229810: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=96;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd229811: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=15;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd229812: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=34;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd229813: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=6;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd229814: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=60;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd229815: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd229957: begin  
rid<=1;
end
19'd229958: begin  
end
19'd229959: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd229960: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd229961: begin  
rid<=0;
end
19'd230101: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=90;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=23822;
 end   
19'd230102: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=76;
   mapp<=59;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=31179;
 end   
19'd230103: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=94;
   mapp<=13;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=30001;
 end   
19'd230104: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=81;
   mapp<=70;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=36928;
 end   
19'd230105: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=92;
   mapp<=71;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=37889;
 end   
19'd230106: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=46;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd230107: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=64;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd230108: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd230109: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd230110: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd230111: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd230112: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=76;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=41510;
 end   
19'd230113: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=65;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=49573;
 end   
19'd230114: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=39;
   mapp<=61;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=44474;
 end   
19'd230115: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=7;
   mapp<=60;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=53538;
 end   
19'd230116: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=34;
   mapp<=12;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=53760;
 end   
19'd230117: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=13;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd230118: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=74;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd230119: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd230120: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd230121: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd230122: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd230123: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd230265: begin  
rid<=1;
end
19'd230266: begin  
end
19'd230267: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd230268: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd230269: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd230270: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd230271: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd230272: begin  
rid<=0;
end
19'd230401: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=93;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7953;
 end   
19'd230402: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=18;
   mapp<=47;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12039;
 end   
19'd230403: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=68;
   mapp<=31;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11035;
 end   
19'd230404: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=62;
   mapp<=62;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=15256;
 end   
19'd230405: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=36;
   mapp<=14;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=11594;
 end   
19'd230406: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=56;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=13790;
 end   
19'd230407: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd230408: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd230409: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd230410: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd230411: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=58;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=24990;
 end   
19'd230412: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=69;
   mapp<=58;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=25275;
 end   
19'd230413: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=96;
   mapp<=71;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=24531;
 end   
19'd230414: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=7;
   mapp<=4;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=29654;
 end   
19'd230415: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=45;
   mapp<=77;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=26066;
 end   
19'd230416: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=90;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=24593;
 end   
19'd230417: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd230418: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd230419: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd230420: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd230421: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd230563: begin  
rid<=1;
end
19'd230564: begin  
end
19'd230565: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd230566: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd230567: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd230568: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd230569: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd230570: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd230571: begin  
rid<=0;
end
19'd230701: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=17;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5131;
 end   
19'd230702: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=23;
   mapp<=54;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7925;
 end   
19'd230703: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=50;
   mapp<=72;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8952;
 end   
19'd230704: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=67;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd230705: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd230706: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=53;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=21768;
 end   
19'd230707: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=84;
   mapp<=80;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=24473;
 end   
19'd230708: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=63;
   mapp<=96;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=18895;
 end   
19'd230709: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=56;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd230710: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=9;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd230711: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd230853: begin  
rid<=1;
end
19'd230854: begin  
end
19'd230855: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd230856: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd230857: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd230858: begin  
rid<=0;
end
19'd231001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=39;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3366;
 end   
19'd231002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=40;
   mapp<=51;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2559;
 end   
19'd231003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=14;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1446;
 end   
19'd231004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=22;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=2248;
 end   
19'd231005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd231006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=54;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=4558;
 end   
19'd231007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=28;
   mapp<=31;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=5997;
 end   
19'd231008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=63;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=5604;
 end   
19'd231009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=27;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=3762;
 end   
19'd231010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd231011: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd231153: begin  
rid<=1;
end
19'd231154: begin  
end
19'd231155: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd231156: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd231157: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd231158: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd231159: begin  
rid<=0;
end
19'd231301: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=36;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13057;
 end   
19'd231302: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=92;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=14196;
 end   
19'd231303: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=91;
   mapp<=23;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12798;
 end   
19'd231304: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=64;
   mapp<=66;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=13411;
 end   
19'd231305: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=19;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd231306: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=31;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd231307: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=98;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd231308: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=19;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=24295;
 end   
19'd231309: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=38;
   mapp<=39;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=24336;
 end   
19'd231310: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=21;
   mapp<=50;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=24983;
 end   
19'd231311: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=93;
   mapp<=93;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=22013;
 end   
19'd231312: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=49;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd231313: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=65;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd231314: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd231315: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd231457: begin  
rid<=1;
end
19'd231458: begin  
end
19'd231459: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd231460: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd231461: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd231462: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd231463: begin  
rid<=0;
end
19'd231601: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=80;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=27292;
 end   
19'd231602: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=1;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=21565;
 end   
19'd231603: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=71;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd231604: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=39;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd231605: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=53;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd231606: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=29;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd231607: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=56;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd231608: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=59;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd231609: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=73;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd231610: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd231611: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=91;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=59090;
 end   
19'd231612: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=15;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=56000;
 end   
19'd231613: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=84;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd231614: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=72;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd231615: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=37;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd231616: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=84;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd231617: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=32;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd231618: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=12;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd231619: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=71;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd231620: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd231621: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd231763: begin  
rid<=1;
end
19'd231764: begin  
end
19'd231765: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd231766: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd231767: begin  
rid<=0;
end
19'd231901: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=72;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12321;
 end   
19'd231902: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=91;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10779;
 end   
19'd231903: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=52;
   mapp<=44;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10512;
 end   
19'd231904: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=20;
   mapp<=34;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=14913;
 end   
19'd231905: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=97;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=14181;
 end   
19'd231906: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=96;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd231907: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd231908: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=30;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd231909: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=48;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=22069;
 end   
19'd231910: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=38;
   mapp<=38;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=17560;
 end   
19'd231911: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=63;
   mapp<=47;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15684;
 end   
19'd231912: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=43;
   mapp<=93;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=21770;
 end   
19'd231913: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=14;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=20773;
 end   
19'd231914: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd231915: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=49;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd231916: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd231917: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd232059: begin  
rid<=1;
end
19'd232060: begin  
end
19'd232061: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd232062: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd232063: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd232064: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd232065: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd232066: begin  
rid<=0;
end
19'd232201: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=16;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14986;
 end   
19'd232202: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=42;
   mapp<=49;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=13314;
 end   
19'd232203: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=52;
   mapp<=0;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=19917;
 end   
19'd232204: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=35;
   mapp<=61;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=11491;
 end   
19'd232205: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=20;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd232206: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=41;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd232207: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=25;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd232208: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=84;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd232209: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=33;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd232210: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=69;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd232211: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=28;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd232212: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=70;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=30490;
 end   
19'd232213: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=1;
   mapp<=70;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=30206;
 end   
19'd232214: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=99;
   mapp<=40;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=37522;
 end   
19'd232215: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=43;
   mapp<=68;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=27844;
 end   
19'd232216: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=18;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd232217: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=28;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd232218: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=9;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd232219: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=55;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd232220: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=17;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd232221: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=64;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd232222: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=68;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd232223: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd232365: begin  
rid<=1;
end
19'd232366: begin  
end
19'd232367: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd232368: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd232369: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd232370: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd232371: begin  
rid<=0;
end
19'd232501: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=46;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2830;
 end   
19'd232502: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=15;
   mapp<=20;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=975;
 end   
19'd232503: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=3;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1553;
 end   
19'd232504: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=93;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5103;
 end   
19'd232505: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=53;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2703;
 end   
19'd232506: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=15;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=1055;
 end   
19'd232507: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=21;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=1656;
 end   
19'd232508: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd232509: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=16;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=6778;
 end   
19'd232510: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=34;
   mapp<=78;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=5113;
 end   
19'd232511: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=85;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=5157;
 end   
19'd232512: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=66;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6703;
 end   
19'd232513: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=16;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=4727;
 end   
19'd232514: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=52;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=5185;
 end   
19'd232515: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=97;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=5384;
 end   
19'd232516: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd232517: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd232659: begin  
rid<=1;
end
19'd232660: begin  
end
19'd232661: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd232662: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd232663: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd232664: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd232665: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd232666: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd232667: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd232668: begin  
rid<=0;
end
19'd232801: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=3;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=19931;
 end   
19'd232802: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=94;
   mapp<=80;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11871;
 end   
19'd232803: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=23;
   mapp<=29;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=15568;
 end   
19'd232804: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=80;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd232805: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=90;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd232806: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=31;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd232807: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=88;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd232808: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=78;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd232809: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd232810: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd232811: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=31;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=44604;
 end   
19'd232812: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=2;
   mapp<=31;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=31762;
 end   
19'd232813: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=94;
   mapp<=95;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=40648;
 end   
19'd232814: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=33;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd232815: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=70;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd232816: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=56;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd232817: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=80;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd232818: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=60;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd232819: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd232820: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd232821: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd232963: begin  
rid<=1;
end
19'd232964: begin  
end
19'd232965: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd232966: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd232967: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd232968: begin  
rid<=0;
end
19'd233101: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=90;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11946;
 end   
19'd233102: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=22;
   mapp<=9;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4176;
 end   
19'd233103: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=68;
   mapp<=51;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10830;
 end   
19'd233104: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=30;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7014;
 end   
19'd233105: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=84;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=13123;
 end   
19'd233106: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=68;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=10305;
 end   
19'd233107: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=93;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=9786;
 end   
19'd233108: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=62;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=8636;
 end   
19'd233109: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=12;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=2588;
 end   
19'd233110: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=54;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd233111: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=18;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd233112: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=60;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=20569;
 end   
19'd233113: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=41;
   mapp<=86;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12843;
 end   
19'd233114: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=69;
   mapp<=53;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=18027;
 end   
19'd233115: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=33;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=16856;
 end   
19'd233116: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=51;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=22551;
 end   
19'd233117: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=88;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=15940;
 end   
19'd233118: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=12;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=15176;
 end   
19'd233119: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=47;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=14399;
 end   
19'd233120: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=20;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=11720;
 end   
19'd233121: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=55;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd233122: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=74;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd233123: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd233265: begin  
rid<=1;
end
19'd233266: begin  
end
19'd233267: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd233268: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd233269: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd233270: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd233271: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd233272: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd233273: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd233274: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd233275: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd233276: begin  
rid<=0;
end
19'd233401: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=32;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6724;
 end   
19'd233402: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=68;
   mapp<=63;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5989;
 end   
19'd233403: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=7;
   mapp<=28;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2694;
 end   
19'd233404: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=12;
   mapp<=1;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4037;
 end   
19'd233405: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=28;
   mapp<=10;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6731;
 end   
19'd233406: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=69;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7434;
 end   
19'd233407: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd233408: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd233409: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd233410: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd233411: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=94;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=18562;
 end   
19'd233412: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=74;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=14236;
 end   
19'd233413: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=81;
   mapp<=28;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=11589;
 end   
19'd233414: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=35;
   mapp<=16;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=17423;
 end   
19'd233415: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=46;
   mapp<=21;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=18338;
 end   
19'd233416: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=86;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=22621;
 end   
19'd233417: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd233418: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd233419: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd233420: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd233421: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd233563: begin  
rid<=1;
end
19'd233564: begin  
end
19'd233565: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd233566: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd233567: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd233568: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd233569: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd233570: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd233571: begin  
rid<=0;
end
19'd233701: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=71;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=26318;
 end   
19'd233702: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=78;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=22740;
 end   
19'd233703: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=0;
   mapp<=87;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=18960;
 end   
19'd233704: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=56;
   mapp<=17;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=22896;
 end   
19'd233705: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=76;
   mapp<=58;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=30067;
 end   
19'd233706: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=80;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd233707: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=98;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd233708: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=36;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd233709: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd233710: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd233711: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=98;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd233712: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=14;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=36109;
 end   
19'd233713: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=37;
   mapp<=49;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=37834;
 end   
19'd233714: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=51;
   mapp<=36;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=40780;
 end   
19'd233715: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=67;
   mapp<=51;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=38810;
 end   
19'd233716: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=32;
   mapp<=33;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=40779;
 end   
19'd233717: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=6;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd233718: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=9;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd233719: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=71;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd233720: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=96;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd233721: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=13;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd233722: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd233723: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd233865: begin  
rid<=1;
end
19'd233866: begin  
end
19'd233867: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd233868: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd233869: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd233870: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd233871: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd233872: begin  
rid<=0;
end
19'd234001: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=43;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2881;
 end   
19'd234002: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=4;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=278;
 end   
19'd234003: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=43;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2901;
 end   
19'd234004: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=92;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6194;
 end   
19'd234005: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=67;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4529;
 end   
19'd234006: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=68;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=4606;
 end   
19'd234007: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=70;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=4750;
 end   
19'd234008: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=2;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=204;
 end   
19'd234009: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=51;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5839;
 end   
19'd234010: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=91;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=5556;
 end   
19'd234011: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=6;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=3249;
 end   
19'd234012: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=33;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=8108;
 end   
19'd234013: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=11;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=5167;
 end   
19'd234014: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=90;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=9826;
 end   
19'd234015: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=79;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=9332;
 end   
19'd234016: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=60;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=3684;
 end   
19'd234017: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd234159: begin  
rid<=1;
end
19'd234160: begin  
end
19'd234161: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd234162: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd234163: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd234164: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd234165: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd234166: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd234167: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd234168: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd234169: begin  
rid<=0;
end
19'd234301: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=84;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=18502;
 end   
19'd234302: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=97;
   mapp<=55;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=22053;
 end   
19'd234303: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=75;
   mapp<=66;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12496;
 end   
19'd234304: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=85;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd234305: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=50;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd234306: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=91;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd234307: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=13;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd234308: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=74;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=36114;
 end   
19'd234309: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=16;
   mapp<=4;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=36165;
 end   
19'd234310: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=45;
   mapp<=84;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=32185;
 end   
19'd234311: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=66;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd234312: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=88;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd234313: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=78;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd234314: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=99;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd234315: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd234457: begin  
rid<=1;
end
19'd234458: begin  
end
19'd234459: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd234460: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd234461: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd234462: begin  
rid<=0;
end
19'd234601: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=60;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=22323;
 end   
19'd234602: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=54;
   mapp<=69;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=24576;
 end   
19'd234603: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=39;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd234604: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=18;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd234605: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=53;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd234606: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=96;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd234607: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=75;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd234608: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=53;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd234609: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=4;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd234610: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd234611: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=77;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=40353;
 end   
19'd234612: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=99;
   mapp<=23;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=39053;
 end   
19'd234613: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=19;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd234614: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=69;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd234615: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=76;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd234616: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=69;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd234617: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=21;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd234618: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=20;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd234619: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd234620: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd234621: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd234763: begin  
rid<=1;
end
19'd234764: begin  
end
19'd234765: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd234766: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd234767: begin  
rid<=0;
end
19'd234901: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=30;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12527;
 end   
19'd234902: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=66;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12860;
 end   
19'd234903: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=83;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd234904: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=3;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd234905: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=42;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=18666;
 end   
19'd234906: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=28;
   mapp<=84;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18383;
 end   
19'd234907: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=35;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd234908: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=35;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd234909: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd235051: begin  
rid<=1;
end
19'd235052: begin  
end
19'd235053: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd235054: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd235055: begin  
rid<=0;
end
19'd235201: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=75;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7904;
 end   
19'd235202: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=54;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd235203: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=4;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd235204: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=83;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd235205: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=11;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd235206: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=10;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd235207: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=85;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=21517;
 end   
19'd235208: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=24;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd235209: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=20;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd235210: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=59;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd235211: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=24;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd235212: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=79;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd235213: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd235355: begin  
rid<=1;
end
19'd235356: begin  
end
19'd235357: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd235358: begin  
rid<=0;
end
19'd235501: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=73;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=24725;
 end   
19'd235502: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=12;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd235503: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=83;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd235504: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=76;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd235505: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=69;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd235506: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=78;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd235507: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=23;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd235508: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=36;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd235509: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=36;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd235510: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=77;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd235511: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=55;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=43001;
 end   
19'd235512: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=50;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd235513: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=66;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd235514: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=17;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd235515: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=4;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd235516: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=43;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd235517: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=21;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd235518: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=33;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd235519: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=23;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd235520: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=42;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd235521: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd235663: begin  
rid<=1;
end
19'd235664: begin  
end
19'd235665: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd235666: begin  
rid<=0;
end
19'd235801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=56;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4312;
 end   
19'd235802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=12;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=682;
 end   
19'd235803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=81;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4556;
 end   
19'd235804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=65;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3670;
 end   
19'd235805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=59;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3344;
 end   
19'd235806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=33;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=1898;
 end   
19'd235807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=89;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8406;
 end   
19'd235808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=3797;
 end   
19'd235809: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=95;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=13011;
 end   
19'd235810: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=67;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=9633;
 end   
19'd235811: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=74;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=9930;
 end   
19'd235812: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=89;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=9819;
 end   
19'd235813: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd235955: begin  
rid<=1;
end
19'd235956: begin  
end
19'd235957: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd235958: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd235959: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd235960: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd235961: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd235962: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd235963: begin  
rid<=0;
end
19'd236101: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=24;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6343;
 end   
19'd236102: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=39;
   mapp<=34;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6579;
 end   
19'd236103: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=55;
   mapp<=55;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7312;
 end   
19'd236104: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=16;
   mapp<=16;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=8536;
 end   
19'd236105: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=52;
   mapp<=8;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=10139;
 end   
19'd236106: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=50;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=12478;
 end   
19'd236107: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=79;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=12692;
 end   
19'd236108: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd236109: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd236110: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd236111: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd236112: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=83;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=29440;
 end   
19'd236113: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=84;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=26970;
 end   
19'd236114: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=13;
   mapp<=66;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=28944;
 end   
19'd236115: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=85;
   mapp<=86;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=32959;
 end   
19'd236116: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=63;
   mapp<=98;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=26930;
 end   
19'd236117: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=33;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=27565;
 end   
19'd236118: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=77;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=29634;
 end   
19'd236119: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd236120: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd236121: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd236122: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd236123: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd236265: begin  
rid<=1;
end
19'd236266: begin  
end
19'd236267: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd236268: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd236269: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd236270: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd236271: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd236272: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd236273: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd236274: begin  
rid<=0;
end
19'd236401: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=77;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7084;
 end   
19'd236402: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=96;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7402;
 end   
19'd236403: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=39;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3023;
 end   
19'd236404: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=10;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=800;
 end   
19'd236405: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=13;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1041;
 end   
19'd236406: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=1;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=127;
 end   
19'd236407: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=29;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=9607;
 end   
19'd236408: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=81;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=9751;
 end   
19'd236409: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=93;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=5720;
 end   
19'd236410: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=58;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=2482;
 end   
19'd236411: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=97;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=3854;
 end   
19'd236412: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=10;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=417;
 end   
19'd236413: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd236555: begin  
rid<=1;
end
19'd236556: begin  
end
19'd236557: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd236558: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd236559: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd236560: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd236561: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd236562: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd236563: begin  
rid<=0;
end
19'd236701: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=42;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13070;
 end   
19'd236702: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=10;
   mapp<=31;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12430;
 end   
19'd236703: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=6;
   mapp<=38;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=14468;
 end   
19'd236704: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=82;
   mapp<=12;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=18813;
 end   
19'd236705: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=56;
   mapp<=37;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=18189;
 end   
19'd236706: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=56;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd236707: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=40;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd236708: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=66;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd236709: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=36;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd236710: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd236711: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd236712: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=76;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=28493;
 end   
19'd236713: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=56;
   mapp<=23;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=25614;
 end   
19'd236714: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=94;
   mapp<=46;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=25403;
 end   
19'd236715: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=55;
   mapp<=86;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=31488;
 end   
19'd236716: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=72;
   mapp<=29;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=28761;
 end   
19'd236717: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=11;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd236718: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=83;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd236719: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=5;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd236720: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=79;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd236721: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=60;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd236722: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=87;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd236723: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd236865: begin  
rid<=1;
end
19'd236866: begin  
end
19'd236867: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd236868: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd236869: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd236870: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd236871: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd236872: begin  
rid<=0;
end
19'd237001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=85;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6801;
 end   
19'd237002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=96;
   mapp<=51;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8046;
 end   
19'd237003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=92;
   mapp<=8;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6047;
 end   
19'd237004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=10;
   mapp<=59;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4160;
 end   
19'd237005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=12;
   mapp<=27;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=11368;
 end   
19'd237006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=84;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7221;
 end   
19'd237007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=7;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd237008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd237009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=63;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd237010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=79;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd237011: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=42;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=15451;
 end   
19'd237012: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=53;
   mapp<=92;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=17745;
 end   
19'd237013: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=53;
   mapp<=20;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=9822;
 end   
19'd237014: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=5;
   mapp<=88;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=12483;
 end   
19'd237015: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=41;
   mapp<=36;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=16787;
 end   
19'd237016: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=3;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=12774;
 end   
19'd237017: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd237018: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=39;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd237019: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=7;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd237020: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=27;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd237021: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd237163: begin  
rid<=1;
end
19'd237164: begin  
end
19'd237165: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd237166: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd237167: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd237168: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd237169: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd237170: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd237171: begin  
rid<=0;
end
19'd237301: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=90;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7200;
 end   
19'd237302: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=52;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4170;
 end   
19'd237303: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=17;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1380;
 end   
19'd237304: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=88;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7070;
 end   
19'd237305: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=15;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1240;
 end   
19'd237306: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=50;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=4050;
 end   
19'd237307: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=42;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=3420;
 end   
19'd237308: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=27;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=2230;
 end   
19'd237309: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=86;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8490;
 end   
19'd237310: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=49;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=4905;
 end   
19'd237311: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=91;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=2745;
 end   
19'd237312: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=24;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=7430;
 end   
19'd237313: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=32;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=1720;
 end   
19'd237314: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=33;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=4545;
 end   
19'd237315: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=93;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=4815;
 end   
19'd237316: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=74;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=3340;
 end   
19'd237317: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd237459: begin  
rid<=1;
end
19'd237460: begin  
end
19'd237461: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd237462: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd237463: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd237464: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd237465: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd237466: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd237467: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd237468: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd237469: begin  
rid<=0;
end
19'd237601: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=57;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7108;
 end   
19'd237602: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=26;
   mapp<=98;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5030;
 end   
19'd237603: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=30;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10946;
 end   
19'd237604: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=87;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=10812;
 end   
19'd237605: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=39;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3846;
 end   
19'd237606: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=7;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=5216;
 end   
19'd237607: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=47;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=4898;
 end   
19'd237608: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=11;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=10456;
 end   
19'd237609: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=97;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=12838;
 end   
19'd237610: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=51;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd237611: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=36;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=9592;
 end   
19'd237612: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=8;
   mapp<=45;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=9777;
 end   
19'd237613: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=95;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=17091;
 end   
19'd237614: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=12;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=13770;
 end   
19'd237615: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=50;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=7966;
 end   
19'd237616: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=26;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=8730;
 end   
19'd237617: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=44;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=10239;
 end   
19'd237618: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=61;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=17250;
 end   
19'd237619: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=71;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=19907;
 end   
19'd237620: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=64;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd237621: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd237763: begin  
rid<=1;
end
19'd237764: begin  
end
19'd237765: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd237766: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd237767: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd237768: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd237769: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd237770: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd237771: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd237772: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd237773: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd237774: begin  
rid<=0;
end
19'd237901: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=75;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=19666;
 end   
19'd237902: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=68;
   mapp<=99;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=20352;
 end   
19'd237903: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=92;
   mapp<=72;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=14585;
 end   
19'd237904: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=17;
   mapp<=45;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=15421;
 end   
19'd237905: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=62;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd237906: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd237907: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd237908: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd237909: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=57;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=30896;
 end   
19'd237910: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=43;
   mapp<=13;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=28751;
 end   
19'd237911: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=55;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=22756;
 end   
19'd237912: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=44;
   mapp<=53;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=21794;
 end   
19'd237913: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=49;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd237914: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd237915: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd237916: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd237917: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd238059: begin  
rid<=1;
end
19'd238060: begin  
end
19'd238061: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd238062: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd238063: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd238064: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd238065: begin  
rid<=0;
end
19'd238201: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=50;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9895;
 end   
19'd238202: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=37;
   mapp<=65;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10507;
 end   
19'd238203: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=85;
   mapp<=72;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=15642;
 end   
19'd238204: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=54;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd238205: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd238206: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd238207: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=88;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=31715;
 end   
19'd238208: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=96;
   mapp<=53;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=30241;
 end   
19'd238209: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=96;
   mapp<=99;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=34728;
 end   
19'd238210: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=50;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd238211: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd238212: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd238213: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd238355: begin  
rid<=1;
end
19'd238356: begin  
end
19'd238357: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd238358: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd238359: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd238360: begin  
rid<=0;
end
19'd238501: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=76;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4256;
 end   
19'd238502: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=79;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6014;
 end   
19'd238503: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=3;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=248;
 end   
19'd238504: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=44;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3374;
 end   
19'd238505: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=17;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1332;
 end   
19'd238506: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=27;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=4364;
 end   
19'd238507: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8579;
 end   
19'd238508: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=30;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=1058;
 end   
19'd238509: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=74;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=5372;
 end   
19'd238510: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=89;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=3735;
 end   
19'd238511: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd238653: begin  
rid<=1;
end
19'd238654: begin  
end
19'd238655: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd238656: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd238657: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd238658: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd238659: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd238660: begin  
rid<=0;
end
19'd238801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=3;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11967;
 end   
19'd238802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=88;
   mapp<=18;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=17845;
 end   
19'd238803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=44;
   mapp<=21;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=13828;
 end   
19'd238804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=42;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd238805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=89;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd238806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=7;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd238807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd238808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=98;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd238809: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=98;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=38687;
 end   
19'd238810: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=36;
   mapp<=82;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=44951;
 end   
19'd238811: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=67;
   mapp<=91;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=41246;
 end   
19'd238812: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=51;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd238813: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=85;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd238814: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=83;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd238815: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=76;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd238816: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=33;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd238817: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd238959: begin  
rid<=1;
end
19'd238960: begin  
end
19'd238961: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd238962: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd238963: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd238964: begin  
rid<=0;
end
19'd239101: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=70;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8208;
 end   
19'd239102: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=18;
   mapp<=71;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8608;
 end   
19'd239103: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=96;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12932;
 end   
19'd239104: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=48;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6273;
 end   
19'd239105: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=21;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=8935;
 end   
19'd239106: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=96;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=13388;
 end   
19'd239107: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=54;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=9737;
 end   
19'd239108: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=61;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=11505;
 end   
19'd239109: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=76;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd239110: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=91;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14704;
 end   
19'd239111: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=28;
   mapp<=76;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12384;
 end   
19'd239112: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=32;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=16672;
 end   
19'd239113: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=29;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=13213;
 end   
19'd239114: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=73;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=17759;
 end   
19'd239115: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=70;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=23208;
 end   
19'd239116: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=85;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=19137;
 end   
19'd239117: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=70;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=17069;
 end   
19'd239118: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=29;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd239119: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd239261: begin  
rid<=1;
end
19'd239262: begin  
end
19'd239263: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd239264: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd239265: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd239266: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd239267: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd239268: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd239269: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd239270: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd239271: begin  
rid<=0;
end
19'd239401: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=33;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3252;
 end   
19'd239402: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=78;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3122;
 end   
19'd239403: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=70;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2500;
 end   
19'd239404: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=55;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3850;
 end   
19'd239405: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=90;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2000;
 end   
19'd239406: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=40;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=3730;
 end   
19'd239407: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=88;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=4212;
 end   
19'd239408: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=95;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd239409: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=60;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7557;
 end   
19'd239410: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=99;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=5418;
 end   
19'd239411: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=26;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=3774;
 end   
19'd239412: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=26;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=5859;
 end   
19'd239413: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=47;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=5213;
 end   
19'd239414: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=73;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=7587;
 end   
19'd239415: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=81;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=7621;
 end   
19'd239416: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=65;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd239417: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd239559: begin  
rid<=1;
end
19'd239560: begin  
end
19'd239561: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd239562: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd239563: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd239564: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd239565: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd239566: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd239567: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd239568: begin  
rid<=0;
end
19'd239701: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=33;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7920;
 end   
19'd239702: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=93;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6271;
 end   
19'd239703: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=40;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9245;
 end   
19'd239704: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd239705: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=65;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17335;
 end   
19'd239706: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=55;
   mapp<=66;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=15731;
 end   
19'd239707: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=94;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=17390;
 end   
19'd239708: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd239709: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd239851: begin  
rid<=1;
end
19'd239852: begin  
end
19'd239853: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd239854: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd239855: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd239856: begin  
rid<=0;
end
19'd240001: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=13;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8820;
 end   
19'd240002: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=76;
   mapp<=16;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12136;
 end   
19'd240003: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=11;
   mapp<=41;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10250;
 end   
19'd240004: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=67;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd240005: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=76;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd240006: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=37;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd240007: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=53;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd240008: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=42;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd240009: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=88;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=20624;
 end   
19'd240010: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=29;
   mapp<=33;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=24927;
 end   
19'd240011: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=12;
   mapp<=59;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=24429;
 end   
19'd240012: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=73;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd240013: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=94;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd240014: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=84;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd240015: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=59;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd240016: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=74;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd240017: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd240159: begin  
rid<=1;
end
19'd240160: begin  
end
19'd240161: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd240162: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd240163: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd240164: begin  
rid<=0;
end
19'd240301: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=60;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8675;
 end   
19'd240302: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=42;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6820;
 end   
19'd240303: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=31;
   mapp<=11;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9056;
 end   
19'd240304: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=79;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=13748;
 end   
19'd240305: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=81;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd240306: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=93;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd240307: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=38;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14508;
 end   
19'd240308: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=50;
   mapp<=60;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=13045;
 end   
19'd240309: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=37;
   mapp<=17;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15459;
 end   
19'd240310: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=65;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=19305;
 end   
19'd240311: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=21;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd240312: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=31;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd240313: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd240455: begin  
rid<=1;
end
19'd240456: begin  
end
19'd240457: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd240458: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd240459: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd240460: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd240461: begin  
rid<=0;
end
19'd240601: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=23;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5304;
 end   
19'd240602: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=76;
   mapp<=26;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9197;
 end   
19'd240603: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=25;
   mapp<=74;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8420;
 end   
19'd240604: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=26;
   mapp<=25;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=9921;
 end   
19'd240605: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=90;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=10389;
 end   
19'd240606: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=98;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=3285;
 end   
19'd240607: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=1;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=4358;
 end   
19'd240608: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd240609: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd240610: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd240611: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=18;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16643;
 end   
19'd240612: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=76;
   mapp<=28;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=17776;
 end   
19'd240613: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=89;
   mapp<=27;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=22614;
 end   
19'd240614: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=94;
   mapp<=55;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=25849;
 end   
19'd240615: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=12;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=29909;
 end   
19'd240616: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=90;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=21723;
 end   
19'd240617: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=64;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=23283;
 end   
19'd240618: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd240619: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd240620: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd240621: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd240763: begin  
rid<=1;
end
19'd240764: begin  
end
19'd240765: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd240766: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd240767: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd240768: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd240769: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd240770: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd240771: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd240772: begin  
rid<=0;
end
19'd240901: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=87;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7917;
 end   
19'd240902: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=0;
   mapp<=92;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8014;
 end   
19'd240903: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=17;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8699;
 end   
19'd240904: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=0;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=9595;
 end   
19'd240905: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd241047: begin  
rid<=1;
end
19'd241048: begin  
end
19'd241049: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd241050: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd241051: begin  
rid<=0;
end
19'd241201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=45;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5023;
 end   
19'd241202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=38;
   mapp<=18;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11038;
 end   
19'd241203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=13;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd241204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=92;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd241205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=98;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14443;
 end   
19'd241206: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=77;
   mapp<=18;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=19891;
 end   
19'd241207: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=74;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd241208: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=71;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd241209: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd241351: begin  
rid<=1;
end
19'd241352: begin  
end
19'd241353: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd241354: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd241355: begin  
rid<=0;
end
19'd241501: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=17;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2187;
 end   
19'd241502: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=1;
   mapp<=70;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7206;
 end   
19'd241503: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=26;
   mapp<=22;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4336;
 end   
19'd241504: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=87;
   mapp<=16;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=8263;
 end   
19'd241505: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=64;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=10185;
 end   
19'd241506: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=26;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6109;
 end   
19'd241507: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=83;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=9811;
 end   
19'd241508: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=79;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=9962;
 end   
19'd241509: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd241510: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd241511: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd241512: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=28;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8710;
 end   
19'd241513: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=39;
   mapp<=39;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=16077;
 end   
19'd241514: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=34;
   mapp<=23;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=10000;
 end   
19'd241515: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=69;
   mapp<=36;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=17638;
 end   
19'd241516: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=82;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=17779;
 end   
19'd241517: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=12;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=16570;
 end   
19'd241518: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=69;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=19933;
 end   
19'd241519: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=36;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=18455;
 end   
19'd241520: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd241521: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd241522: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd241523: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd241665: begin  
rid<=1;
end
19'd241666: begin  
end
19'd241667: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd241668: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd241669: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd241670: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd241671: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd241672: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd241673: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd241674: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd241675: begin  
rid<=0;
end
19'd241801: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=1;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14750;
 end   
19'd241802: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=72;
   mapp<=31;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15670;
 end   
19'd241803: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=82;
   mapp<=95;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11987;
 end   
19'd241804: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=22;
   mapp<=29;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=13351;
 end   
19'd241805: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=40;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd241806: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=45;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd241807: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=57;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd241808: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd241809: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd241810: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd241811: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=73;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=29740;
 end   
19'd241812: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=59;
   mapp<=8;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=32169;
 end   
19'd241813: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=46;
   mapp<=86;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=29347;
 end   
19'd241814: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=77;
   mapp<=25;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=29569;
 end   
19'd241815: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=15;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd241816: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=11;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd241817: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=80;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd241818: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd241819: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd241820: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd241821: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd241963: begin  
rid<=1;
end
19'd241964: begin  
end
19'd241965: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd241966: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd241967: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd241968: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd241969: begin  
rid<=0;
end
19'd242101: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=2;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2906;
 end   
19'd242102: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=58;
   mapp<=31;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3716;
 end   
19'd242103: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=14;
   mapp<=74;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1538;
 end   
19'd242104: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=16;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=2081;
 end   
19'd242105: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=7;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2743;
 end   
19'd242106: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=17;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=8720;
 end   
19'd242107: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=26;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=5810;
 end   
19'd242108: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=98;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd242109: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=24;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd242110: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=82;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14751;
 end   
19'd242111: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=85;
   mapp<=57;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=11573;
 end   
19'd242112: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=6;
   mapp<=5;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=5659;
 end   
19'd242113: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=58;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=10598;
 end   
19'd242114: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=61;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=9382;
 end   
19'd242115: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=22;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=13055;
 end   
19'd242116: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=40;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=11474;
 end   
19'd242117: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd242118: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=31;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd242119: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd242261: begin  
rid<=1;
end
19'd242262: begin  
end
19'd242263: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd242264: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd242265: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd242266: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd242267: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd242268: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd242269: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd242270: begin  
rid<=0;
end
19'd242401: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=97;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16542;
 end   
19'd242402: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=81;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd242403: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=76;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd242404: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=72;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd242405: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=85;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd242406: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=74;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=39961;
 end   
19'd242407: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=80;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd242408: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=72;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd242409: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=96;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd242410: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=1;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd242411: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd242553: begin  
rid<=1;
end
19'd242554: begin  
end
19'd242555: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd242556: begin  
rid<=0;
end
19'd242701: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=11;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13072;
 end   
19'd242702: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=28;
   mapp<=43;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=14089;
 end   
19'd242703: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=37;
   mapp<=52;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11940;
 end   
19'd242704: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=32;
   mapp<=21;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=15719;
 end   
19'd242705: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=58;
   mapp<=70;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=17739;
 end   
19'd242706: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=84;
   mapp<=50;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=16834;
 end   
19'd242707: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd242708: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=15;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd242709: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=87;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd242710: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd242711: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=77;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd242712: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=3;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=26806;
 end   
19'd242713: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=38;
   mapp<=11;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=29462;
 end   
19'd242714: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=51;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=28832;
 end   
19'd242715: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=53;
   mapp<=41;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=34192;
 end   
19'd242716: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=5;
   mapp<=89;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=27560;
 end   
19'd242717: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=73;
   mapp<=96;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=29123;
 end   
19'd242718: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=30;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd242719: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=86;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd242720: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=24;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd242721: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=11;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd242722: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=11;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd242723: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd242865: begin  
rid<=1;
end
19'd242866: begin  
end
19'd242867: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd242868: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd242869: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd242870: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd242871: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd242872: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd242873: begin  
rid<=0;
end
19'd243001: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=94;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13715;
 end   
19'd243002: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=78;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd243003: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=33;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd243004: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=58;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd243005: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=53;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=24809;
 end   
19'd243006: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=93;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd243007: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=25;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd243008: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=54;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd243009: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd243151: begin  
rid<=1;
end
19'd243152: begin  
end
19'd243153: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd243154: begin  
rid<=0;
end
19'd243301: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=13;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=19045;
 end   
19'd243302: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=80;
   mapp<=36;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=19802;
 end   
19'd243303: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=50;
   mapp<=57;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=21483;
 end   
19'd243304: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=46;
   mapp<=91;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=20836;
 end   
19'd243305: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=34;
   mapp<=42;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=18636;
 end   
19'd243306: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=93;
   mapp<=74;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=24779;
 end   
19'd243307: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=45;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd243308: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=59;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd243309: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=65;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd243310: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=33;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd243311: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd243312: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=61;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=36854;
 end   
19'd243313: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=36;
   mapp<=24;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=35569;
 end   
19'd243314: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=64;
   mapp<=43;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=38663;
 end   
19'd243315: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=96;
   mapp<=67;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=38820;
 end   
19'd243316: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=29;
   mapp<=33;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=31839;
 end   
19'd243317: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=96;
   mapp<=48;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=41599;
 end   
19'd243318: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=77;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd243319: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=49;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd243320: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=61;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd243321: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=26;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd243322: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=93;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd243323: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd243465: begin  
rid<=1;
end
19'd243466: begin  
end
19'd243467: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd243468: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd243469: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd243470: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd243471: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd243472: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd243473: begin  
rid<=0;
end
19'd243601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=50;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13250;
 end   
19'd243602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=26;
   mapp<=43;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=14167;
 end   
19'd243603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=73;
   mapp<=54;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12833;
 end   
19'd243604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=40;
   mapp<=91;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=11263;
 end   
19'd243605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=99;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=14615;
 end   
19'd243606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=13;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=9658;
 end   
19'd243607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd243608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd243609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd243610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=58;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=26449;
 end   
19'd243611: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=23;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=22473;
 end   
19'd243612: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=97;
   mapp<=69;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=21443;
 end   
19'd243613: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=18;
   mapp<=65;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=21755;
 end   
19'd243614: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=23;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=25376;
 end   
19'd243615: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=49;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=18942;
 end   
19'd243616: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd243617: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd243618: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd243619: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd243761: begin  
rid<=1;
end
19'd243762: begin  
end
19'd243763: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd243764: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd243765: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd243766: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd243767: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd243768: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd243769: begin  
rid<=0;
end
19'd243901: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6800;
 end   
19'd243902: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=80;
   mapp<=85;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5610;
 end   
19'd243903: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3220;
 end   
19'd243904: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=40;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7710;
 end   
19'd243905: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=96;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1160;
 end   
19'd243906: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=14;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=4050;
 end   
19'd243907: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd243908: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=45;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17285;
 end   
19'd243909: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=75;
   mapp<=96;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=15780;
 end   
19'd243910: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=78;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=7105;
 end   
19'd243911: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=5;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=10260;
 end   
19'd243912: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=31;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=8855;
 end   
19'd243913: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=84;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=12630;
 end   
19'd243914: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd243915: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd244057: begin  
rid<=1;
end
19'd244058: begin  
end
19'd244059: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd244060: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd244061: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd244062: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd244063: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd244064: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd244065: begin  
rid<=0;
end
19'd244201: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=83;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14017;
 end   
19'd244202: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=95;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd244203: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=84;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd244204: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=30;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd244205: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=31;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd244206: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=97;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd244207: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=29;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=37234;
 end   
19'd244208: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=73;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd244209: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=46;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd244210: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=67;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd244211: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=92;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd244212: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=94;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd244213: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd244355: begin  
rid<=1;
end
19'd244356: begin  
end
19'd244357: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd244358: begin  
rid<=0;
end
19'd244501: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=55;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4950;
 end   
19'd244502: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=74;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4080;
 end   
19'd244503: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3870;
 end   
19'd244504: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=50;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=2780;
 end   
19'd244505: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=73;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7578;
 end   
19'd244506: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=64;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8752;
 end   
19'd244507: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=51;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=7593;
 end   
19'd244508: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=20;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=4240;
 end   
19'd244509: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd244651: begin  
rid<=1;
end
19'd244652: begin  
end
19'd244653: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd244654: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd244655: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd244656: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd244657: begin  
rid<=0;
end
19'd244801: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=67;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8944;
 end   
19'd244802: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=18;
   mapp<=85;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10356;
 end   
19'd244803: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=85;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd244804: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=25;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd244805: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=70;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd244806: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=25;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd244807: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=40;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=13865;
 end   
19'd244808: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=48;
   mapp<=33;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=14898;
 end   
19'd244809: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=56;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd244810: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=30;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd244811: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=77;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd244812: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=31;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd244813: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd244955: begin  
rid<=1;
end
19'd244956: begin  
end
19'd244957: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd244958: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd244959: begin  
rid<=0;
end
19'd245101: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=45;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2919;
 end   
19'd245102: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=11;
   mapp<=6;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5385;
 end   
19'd245103: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=54;
   mapp<=37;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4640;
 end   
19'd245104: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=87;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7106;
 end   
19'd245105: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=37;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5344;
 end   
19'd245106: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=51;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=3836;
 end   
19'd245107: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=57;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=3449;
 end   
19'd245108: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd245109: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd245110: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=59;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=9382;
 end   
19'd245111: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=85;
   mapp<=13;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12392;
 end   
19'd245112: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=60;
   mapp<=48;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=13532;
 end   
19'd245113: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=36;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=18160;
 end   
19'd245114: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=50;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=17384;
 end   
19'd245115: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=78;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=13783;
 end   
19'd245116: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=41;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=13303;
 end   
19'd245117: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd245118: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd245119: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd245261: begin  
rid<=1;
end
19'd245262: begin  
end
19'd245263: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd245264: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd245265: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd245266: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd245267: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd245268: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd245269: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd245270: begin  
rid<=0;
end
19'd245401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=99;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9021;
 end   
19'd245402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=84;
   mapp<=19;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9283;
 end   
19'd245403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd245404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=50;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=10121;
 end   
19'd245405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=41;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12891;
 end   
19'd245406: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd245407: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd245549: begin  
rid<=1;
end
19'd245550: begin  
end
19'd245551: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd245552: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd245553: begin  
rid<=0;
end
19'd245701: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=47;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5469;
 end   
19'd245702: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=31;
   mapp<=37;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5321;
 end   
19'd245703: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=41;
   mapp<=16;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6864;
 end   
19'd245704: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=86;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7827;
 end   
19'd245705: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=29;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3091;
 end   
19'd245706: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=1;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=3099;
 end   
19'd245707: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=47;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd245708: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=77;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd245709: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=38;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=15143;
 end   
19'd245710: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=36;
   mapp<=65;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=13506;
 end   
19'd245711: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=73;
   mapp<=76;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15210;
 end   
19'd245712: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=23;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=16849;
 end   
19'd245713: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=45;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=10028;
 end   
19'd245714: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=66;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=6884;
 end   
19'd245715: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=7;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd245716: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=3;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd245717: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd245859: begin  
rid<=1;
end
19'd245860: begin  
end
19'd245861: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd245862: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd245863: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd245864: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd245865: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd245866: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd245867: begin  
rid<=0;
end
19'd246001: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=71;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6035;
 end   
19'd246002: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=46;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3920;
 end   
19'd246003: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=66;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5630;
 end   
19'd246004: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=30;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8285;
 end   
19'd246005: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=30;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=6170;
 end   
19'd246006: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=14;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=6680;
 end   
19'd246007: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd246149: begin  
rid<=1;
end
19'd246150: begin  
end
19'd246151: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd246152: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd246153: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd246154: begin  
rid<=0;
end
19'd246301: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=52;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6664;
 end   
19'd246302: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=17;
   mapp<=7;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=14942;
 end   
19'd246303: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=29;
   mapp<=30;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9784;
 end   
19'd246304: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=20;
   mapp<=87;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=15613;
 end   
19'd246305: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=89;
   mapp<=30;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=10731;
 end   
19'd246306: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=9;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd246307: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=77;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd246308: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=46;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd246309: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=83;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd246310: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=11;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd246311: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=24;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17328;
 end   
19'd246312: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=80;
   mapp<=66;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=26453;
 end   
19'd246313: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=30;
   mapp<=97;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=19376;
 end   
19'd246314: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=7;
   mapp<=70;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=23407;
 end   
19'd246315: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=64;
   mapp<=10;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=19160;
 end   
19'd246316: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=12;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd246317: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=21;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd246318: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=31;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd246319: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd246320: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd246321: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd246463: begin  
rid<=1;
end
19'd246464: begin  
end
19'd246465: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd246466: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd246467: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd246468: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd246469: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd246470: begin  
rid<=0;
end
19'd246601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=10;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5156;
 end   
19'd246602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=87;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9103;
 end   
19'd246603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=99;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8318;
 end   
19'd246604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=84;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4872;
 end   
19'd246605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=46;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6677;
 end   
19'd246606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=71;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=3370;
 end   
19'd246607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=30;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=8103;
 end   
19'd246608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=89;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=6615;
 end   
19'd246609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd246610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=87;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=15092;
 end   
19'd246611: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=33;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18607;
 end   
19'd246612: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=85;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=18056;
 end   
19'd246613: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=71;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=11478;
 end   
19'd246614: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=13;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=8237;
 end   
19'd246615: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=13;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=4864;
 end   
19'd246616: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=11;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=12294;
 end   
19'd246617: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=98;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=17682;
 end   
19'd246618: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd246619: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd246761: begin  
rid<=1;
end
19'd246762: begin  
end
19'd246763: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd246764: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd246765: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd246766: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd246767: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd246768: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd246769: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd246770: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd246771: begin  
rid<=0;
end
19'd246901: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=19;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=642;
 end   
19'd246902: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=2;
   mapp<=55;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2596;
 end   
19'd246903: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=46;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6203;
 end   
19'd246904: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd246905: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=43;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7303;
 end   
19'd246906: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=55;
   mapp<=57;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=10298;
 end   
19'd246907: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=56;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15013;
 end   
19'd246908: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=74;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd246909: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd247051: begin  
rid<=1;
end
19'd247052: begin  
end
19'd247053: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd247054: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd247055: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd247056: begin  
rid<=0;
end
19'd247201: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=29;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16438;
 end   
19'd247202: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=6;
   mapp<=94;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=16611;
 end   
19'd247203: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=62;
   mapp<=92;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=15358;
 end   
19'd247204: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=62;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd247205: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=26;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd247206: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=53;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd247207: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=73;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd247208: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd247209: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd247210: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=96;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=33109;
 end   
19'd247211: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=63;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=36149;
 end   
19'd247212: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=13;
   mapp<=93;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=37376;
 end   
19'd247213: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=13;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd247214: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=38;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd247215: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=27;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd247216: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=37;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd247217: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd247218: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd247219: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd247361: begin  
rid<=1;
end
19'd247362: begin  
end
19'd247363: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd247364: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd247365: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd247366: begin  
rid<=0;
end
19'd247501: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=42;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9583;
 end   
19'd247502: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=67;
   mapp<=71;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10380;
 end   
19'd247503: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=19;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd247504: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=50;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd247505: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=64;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd247506: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd247507: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=9;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=29477;
 end   
19'd247508: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=59;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=33457;
 end   
19'd247509: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=94;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd247510: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=82;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd247511: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=68;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd247512: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=61;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd247513: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd247655: begin  
rid<=1;
end
19'd247656: begin  
end
19'd247657: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd247658: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd247659: begin  
rid<=0;
end
19'd247801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=95;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=446;
 end   
19'd247802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=2;
   mapp<=33;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1800;
 end   
19'd247803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=54;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=797;
 end   
19'd247804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=17;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=263;
 end   
19'd247805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=5;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd247806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=58;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5579;
 end   
19'd247807: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=87;
   mapp<=43;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=6769;
 end   
19'd247808: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=67;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=6361;
 end   
19'd247809: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=92;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=5051;
 end   
19'd247810: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=60;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd247811: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd247953: begin  
rid<=1;
end
19'd247954: begin  
end
19'd247955: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd247956: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd247957: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd247958: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd247959: begin  
rid<=0;
end
19'd248101: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=87;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8609;
 end   
19'd248102: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=15;
   mapp<=1;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=938;
 end   
19'd248103: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=79;
   mapp<=35;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4073;
 end   
19'd248104: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=4;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3718;
 end   
19'd248105: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=12;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=9347;
 end   
19'd248106: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=40;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=9409;
 end   
19'd248107: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=97;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=10050;
 end   
19'd248108: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd248109: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd248110: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=45;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=13245;
 end   
19'd248111: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=52;
   mapp<=4;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=4369;
 end   
19'd248112: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=9;
   mapp<=62;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=7658;
 end   
19'd248113: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=3;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=8157;
 end   
19'd248114: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=71;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=16078;
 end   
19'd248115: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=68;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=12658;
 end   
19'd248116: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=11754;
 end   
19'd248117: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd248118: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd248119: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd248261: begin  
rid<=1;
end
19'd248262: begin  
end
19'd248263: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd248264: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd248265: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd248266: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd248267: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd248268: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd248269: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd248270: begin  
rid<=0;
end
19'd248401: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=62;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2422;
 end   
19'd248402: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=37;
   mapp<=42;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4350;
 end   
19'd248403: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=91;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2722;
 end   
19'd248404: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd248405: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=12;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7114;
 end   
19'd248406: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=77;
   mapp<=60;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8052;
 end   
19'd248407: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=54;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=7306;
 end   
19'd248408: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=71;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd248409: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd248551: begin  
rid<=1;
end
19'd248552: begin  
end
19'd248553: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd248554: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd248555: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd248556: begin  
rid<=0;
end
19'd248701: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=95;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4943;
 end   
19'd248702: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=6;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2080;
 end   
19'd248703: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=37;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2793;
 end   
19'd248704: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=20;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=2594;
 end   
19'd248705: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=33;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3913;
 end   
19'd248706: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=47;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6385;
 end   
19'd248707: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=84;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=4608;
 end   
19'd248708: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=9;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=2575;
 end   
19'd248709: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=43;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=6171;
 end   
19'd248710: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=83;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=8765;
 end   
19'd248711: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=96;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd248712: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=87;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14134;
 end   
19'd248713: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=16;
   mapp<=47;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=7862;
 end   
19'd248714: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=90;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=12416;
 end   
19'd248715: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=19;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=8291;
 end   
19'd248716: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=82;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=14875;
 end   
19'd248717: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=64;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=16447;
 end   
19'd248718: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=82;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=13549;
 end   
19'd248719: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=21;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=8513;
 end   
19'd248720: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=83;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=17183;
 end   
19'd248721: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=63;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=16662;
 end   
19'd248722: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd248723: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd248865: begin  
rid<=1;
end
19'd248866: begin  
end
19'd248867: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd248868: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd248869: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd248870: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd248871: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd248872: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd248873: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd248874: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd248875: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd248876: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd248877: begin  
rid<=0;
end
19'd249001: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=69;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4347;
 end   
19'd249002: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6703;
 end   
19'd249003: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4850;
 end   
19'd249004: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=40;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=2790;
 end   
19'd249005: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=40;
 end   
19'd249006: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=10;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=740;
 end   
19'd249007: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=16;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=1164;
 end   
19'd249008: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=41;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7955;
 end   
19'd249009: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=10680;
 end   
19'd249010: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=55;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=7105;
 end   
19'd249011: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=18;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=3528;
 end   
19'd249012: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=51;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=2131;
 end   
19'd249013: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=61;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=3241;
 end   
19'd249014: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=45;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=3009;
 end   
19'd249015: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd249157: begin  
rid<=1;
end
19'd249158: begin  
end
19'd249159: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd249160: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd249161: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd249162: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd249163: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd249164: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd249165: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd249166: begin  
rid<=0;
end
19'd249301: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=66;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11705;
 end   
19'd249302: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=57;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8845;
 end   
19'd249303: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=21;
   mapp<=23;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11502;
 end   
19'd249304: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=58;
   mapp<=7;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=9404;
 end   
19'd249305: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=74;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd249306: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=19;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd249307: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=65;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd249308: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd249309: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=83;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd249310: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=11;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd249311: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=76;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=32062;
 end   
19'd249312: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=90;
   mapp<=60;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=24982;
 end   
19'd249313: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=16;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=21043;
 end   
19'd249314: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=28;
   mapp<=40;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=20629;
 end   
19'd249315: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=76;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd249316: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=81;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd249317: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=57;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd249318: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=35;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd249319: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=7;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd249320: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=5;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd249321: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd249463: begin  
rid<=1;
end
19'd249464: begin  
end
19'd249465: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd249466: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd249467: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd249468: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd249469: begin  
rid<=0;
end
19'd249601: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=47;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4923;
 end   
19'd249602: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=45;
   mapp<=62;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5941;
 end   
19'd249603: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=70;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd249604: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=26;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd249605: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=48;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8111;
 end   
19'd249606: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=48;
   mapp<=21;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=9662;
 end   
19'd249607: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=1;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd249608: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=77;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd249609: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd249751: begin  
rid<=1;
end
19'd249752: begin  
end
19'd249753: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd249754: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd249755: begin  
rid<=0;
end
19'd249901: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=25;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1875;
 end   
19'd249902: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=36;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=910;
 end   
19'd249903: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=10;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=270;
 end   
19'd249904: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=25;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=655;
 end   
19'd249905: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=9;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=265;
 end   
19'd249906: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=93;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=6153;
 end   
19'd249907: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=9559;
 end   
19'd249908: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=83;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=7989;
 end   
19'd249909: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=88;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=8839;
 end   
19'd249910: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=94;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=9007;
 end   
19'd249911: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd250053: begin  
rid<=1;
end
19'd250054: begin  
end
19'd250055: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd250056: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd250057: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd250058: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd250059: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd250060: begin  
rid<=0;
end
19'd250201: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=61;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10857;
 end   
19'd250202: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=2;
   mapp<=27;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3234;
 end   
19'd250203: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=7;
   mapp<=82;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9794;
 end   
19'd250204: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=70;
   mapp<=77;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=12958;
 end   
19'd250205: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=66;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd250206: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd250207: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd250208: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd250209: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=39;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=21220;
 end   
19'd250210: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=93;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=16931;
 end   
19'd250211: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=62;
   mapp<=56;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=21087;
 end   
19'd250212: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=91;
   mapp<=6;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=32042;
 end   
19'd250213: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=45;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd250214: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd250215: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd250216: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd250217: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd250359: begin  
rid<=1;
end
19'd250360: begin  
end
19'd250361: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd250362: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd250363: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd250364: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd250365: begin  
rid<=0;
end
19'd250501: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=80;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11896;
 end   
19'd250502: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=88;
   mapp<=87;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12417;
 end   
19'd250503: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=89;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5868;
 end   
19'd250504: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=13;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1067;
 end   
19'd250505: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=4;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1731;
 end   
19'd250506: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=17;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=8694;
 end   
19'd250507: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=89;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=6952;
 end   
19'd250508: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=25;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=7572;
 end   
19'd250509: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=71;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd250510: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=74;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17904;
 end   
19'd250511: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=62;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=17366;
 end   
19'd250512: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=35;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=8713;
 end   
19'd250513: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=30;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=3767;
 end   
19'd250514: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=78;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=8222;
 end   
19'd250515: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=97;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=16173;
 end   
19'd250516: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=2;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=7171;
 end   
19'd250517: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=13;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=8643;
 end   
19'd250518: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=14;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd250519: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd250661: begin  
rid<=1;
end
19'd250662: begin  
end
19'd250663: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd250664: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd250665: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd250666: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd250667: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd250668: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd250669: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd250670: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd250671: begin  
rid<=0;
end
19'd250801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=60;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9672;
 end   
19'd250802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=92;
   mapp<=51;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10349;
 end   
19'd250803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=53;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8448;
 end   
19'd250804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=79;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=9953;
 end   
19'd250805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=66;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=7558;
 end   
19'd250806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=40;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=3982;
 end   
19'd250807: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd250808: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=54;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=13930;
 end   
19'd250809: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=95;
   mapp<=38;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12591;
 end   
19'd250810: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=29;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=12482;
 end   
19'd250811: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=97;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=12447;
 end   
19'd250812: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=35;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=10562;
 end   
19'd250813: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=68;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=8370;
 end   
19'd250814: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=94;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd250815: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd250957: begin  
rid<=1;
end
19'd250958: begin  
end
19'd250959: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd250960: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd250961: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd250962: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd250963: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd250964: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd250965: begin  
rid<=0;
end
19'd251101: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=2;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6877;
 end   
19'd251102: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=11;
   mapp<=25;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9366;
 end   
19'd251103: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=89;
   mapp<=8;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10684;
 end   
19'd251104: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=68;
   mapp<=63;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=11585;
 end   
19'd251105: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=78;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd251106: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=71;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd251107: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=91;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd251108: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=87;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd251109: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=94;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=21679;
 end   
19'd251110: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=48;
   mapp<=39;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=21212;
 end   
19'd251111: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=81;
   mapp<=89;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=22377;
 end   
19'd251112: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=57;
   mapp<=41;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=23108;
 end   
19'd251113: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=46;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd251114: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=60;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd251115: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=57;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd251116: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=32;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd251117: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd251259: begin  
rid<=1;
end
19'd251260: begin  
end
19'd251261: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd251262: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd251263: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd251264: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd251265: begin  
rid<=0;
end
19'd251401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=3;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=22533;
 end   
19'd251402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=62;
   mapp<=6;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=20524;
 end   
19'd251403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=15;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd251404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=3;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd251405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=25;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd251406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=60;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd251407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=95;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd251408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=20;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd251409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=40;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd251410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=82;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd251411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd251412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=3;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=47055;
 end   
19'd251413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=38;
   mapp<=98;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=46825;
 end   
19'd251414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=7;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd251415: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=72;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd251416: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=68;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd251417: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=33;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd251418: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=71;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd251419: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=96;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd251420: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=70;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd251421: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=13;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd251422: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd251423: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd251565: begin  
rid<=1;
end
19'd251566: begin  
end
19'd251567: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd251568: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd251569: begin  
rid<=0;
end
19'd251701: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=51;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1089;
 end   
19'd251702: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=70;
   mapp<=9;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6139;
 end   
19'd251703: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=81;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8071;
 end   
19'd251704: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=56;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=9116;
 end   
19'd251705: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=89;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5979;
 end   
19'd251706: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=20;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7370;
 end   
19'd251707: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=90;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=8080;
 end   
19'd251708: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=49;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=4109;
 end   
19'd251709: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=22;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=7152;
 end   
19'd251710: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd251711: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=98;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12031;
 end   
19'd251712: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=61;
   mapp<=38;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=10168;
 end   
19'd251713: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=5;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=14356;
 end   
19'd251714: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=95;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=19585;
 end   
19'd251715: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=19;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=8634;
 end   
19'd251716: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=13;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=14378;
 end   
19'd251717: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=94;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=21745;
 end   
19'd251718: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=73;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=13642;
 end   
19'd251719: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=39;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=16586;
 end   
19'd251720: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd251721: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd251863: begin  
rid<=1;
end
19'd251864: begin  
end
19'd251865: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd251866: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd251867: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd251868: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd251869: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd251870: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd251871: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd251872: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd251873: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd251874: begin  
rid<=0;
end
19'd252001: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=69;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8527;
 end   
19'd252002: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=68;
   mapp<=29;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8819;
 end   
19'd252003: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=81;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd252004: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=55;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=13769;
 end   
19'd252005: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=81;
   mapp<=7;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=15844;
 end   
19'd252006: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=20;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd252007: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd252149: begin  
rid<=1;
end
19'd252150: begin  
end
19'd252151: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd252152: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd252153: begin  
rid<=0;
end
19'd252301: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=26;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2852;
 end   
19'd252302: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=32;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2642;
 end   
19'd252303: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd252304: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=92;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=6789;
 end   
19'd252305: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=97;
   mapp<=33;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8879;
 end   
19'd252306: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd252307: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd252449: begin  
rid<=1;
end
19'd252450: begin  
end
19'd252451: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd252452: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd252453: begin  
rid<=0;
end
19'd252601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=77;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7504;
 end   
19'd252602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=4;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6981;
 end   
19'd252603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=11;
   mapp<=57;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4823;
 end   
19'd252604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=32;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3566;
 end   
19'd252605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=26;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3153;
 end   
19'd252606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=88;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7949;
 end   
19'd252607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=69;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=5978;
 end   
19'd252608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd252609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd252610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=1;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=9265;
 end   
19'd252611: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=18;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=10905;
 end   
19'd252612: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=41;
   mapp<=9;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=10019;
 end   
19'd252613: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=90;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=5796;
 end   
19'd252614: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=87;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=4722;
 end   
19'd252615: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=14;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=9036;
 end   
19'd252616: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=30;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=7800;
 end   
19'd252617: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd252618: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd252619: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd252761: begin  
rid<=1;
end
19'd252762: begin  
end
19'd252763: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd252764: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd252765: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd252766: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd252767: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd252768: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd252769: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd252770: begin  
rid<=0;
end
19'd252901: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=69;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=414;
 end   
19'd252902: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=19;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=433;
 end   
19'd252903: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd253045: begin  
rid<=1;
end
19'd253046: begin  
end
19'd253047: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd253048: begin  
rid<=0;
end
19'd253201: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=54;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3294;
 end   
19'd253202: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=35;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2145;
 end   
19'd253203: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=74;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4534;
 end   
19'd253204: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=24;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1494;
 end   
19'd253205: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=8;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=3814;
 end   
19'd253206: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=12;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=2925;
 end   
19'd253207: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=15;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=5509;
 end   
19'd253208: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=84;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6954;
 end   
19'd253209: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd253351: begin  
rid<=1;
end
19'd253352: begin  
end
19'd253353: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd253354: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd253355: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd253356: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd253357: begin  
rid<=0;
end
19'd253501: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=18;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=15818;
 end   
19'd253502: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=25;
   mapp<=99;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=19561;
 end   
19'd253503: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=97;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd253504: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=67;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd253505: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=3;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd253506: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=3;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd253507: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=60;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd253508: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=1;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd253509: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=59;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=42732;
 end   
19'd253510: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=92;
   mapp<=71;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=42097;
 end   
19'd253511: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=94;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd253512: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=48;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd253513: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=85;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd253514: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=14;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd253515: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=56;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd253516: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=26;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd253517: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd253659: begin  
rid<=1;
end
19'd253660: begin  
end
19'd253661: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd253662: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd253663: begin  
rid<=0;
end
19'd253801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=93;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=34460;
 end   
19'd253802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=87;
   mapp<=98;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=31761;
 end   
19'd253803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=22;
   mapp<=64;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=29351;
 end   
19'd253804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=34;
   mapp<=65;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=31056;
 end   
19'd253805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=91;
   mapp<=63;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=30560;
 end   
19'd253806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=81;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd253807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=59;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd253808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=83;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd253809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd253810: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=35;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd253811: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=39;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd253812: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=14;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=54251;
 end   
19'd253813: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=72;
   mapp<=98;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=63709;
 end   
19'd253814: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=98;
   mapp<=25;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=54375;
 end   
19'd253815: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=21;
   mapp<=74;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=45312;
 end   
19'd253816: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=12;
   mapp<=47;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=55194;
 end   
19'd253817: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=98;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd253818: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=19;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd253819: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=98;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd253820: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=17;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd253821: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=21;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd253822: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=45;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd253823: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd253965: begin  
rid<=1;
end
19'd253966: begin  
end
19'd253967: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd253968: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd253969: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd253970: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd253971: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd253972: begin  
rid<=0;
end
19'd254101: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=25;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3948;
 end   
19'd254102: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=31;
   mapp<=81;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5974;
 end   
19'd254103: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=61;
   mapp<=17;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4408;
 end   
19'd254104: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=31;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5159;
 end   
19'd254105: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=53;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2916;
 end   
19'd254106: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=20;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=3810;
 end   
19'd254107: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=24;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=8745;
 end   
19'd254108: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=88;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=8121;
 end   
19'd254109: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=69;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd254110: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd254111: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=87;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=13569;
 end   
19'd254112: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=79;
   mapp<=57;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=14119;
 end   
19'd254113: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=27;
   mapp<=80;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15159;
 end   
19'd254114: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=49;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=18961;
 end   
19'd254115: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=88;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=13141;
 end   
19'd254116: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=89;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=12215;
 end   
19'd254117: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=27;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=18159;
 end   
19'd254118: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=48;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=15777;
 end   
19'd254119: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=72;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd254120: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=24;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd254121: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd254263: begin  
rid<=1;
end
19'd254264: begin  
end
19'd254265: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd254266: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd254267: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd254268: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd254269: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd254270: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd254271: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd254272: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd254273: begin  
rid<=0;
end
19'd254401: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=51;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10288;
 end   
19'd254402: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=66;
   mapp<=26;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=13273;
 end   
19'd254403: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=38;
   mapp<=96;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8493;
 end   
19'd254404: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=89;
   mapp<=33;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7391;
 end   
19'd254405: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=11;
   mapp<=74;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=9776;
 end   
19'd254406: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=25;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6342;
 end   
19'd254407: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=46;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd254408: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=15;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd254409: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=53;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd254410: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=18;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd254411: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=41;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=28978;
 end   
19'd254412: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=51;
   mapp<=79;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=33234;
 end   
19'd254413: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=95;
   mapp<=30;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=23989;
 end   
19'd254414: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=94;
   mapp<=23;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=27145;
 end   
19'd254415: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=78;
   mapp<=99;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=20723;
 end   
19'd254416: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=55;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=12671;
 end   
19'd254417: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd254418: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=76;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd254419: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd254420: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd254421: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd254563: begin  
rid<=1;
end
19'd254564: begin  
end
19'd254565: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd254566: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd254567: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd254568: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd254569: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd254570: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd254571: begin  
rid<=0;
end
19'd254701: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=91;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9076;
 end   
19'd254702: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=33;
   mapp<=12;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3652;
 end   
19'd254703: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=94;
   mapp<=42;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6900;
 end   
19'd254704: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=19;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4084;
 end   
19'd254705: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=42;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4594;
 end   
19'd254706: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=61;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=4362;
 end   
19'd254707: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=39;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd254708: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd254709: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=13;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12316;
 end   
19'd254710: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=45;
   mapp<=46;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=7724;
 end   
19'd254711: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=6;
   mapp<=26;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=8056;
 end   
19'd254712: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=11;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6278;
 end   
19'd254713: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=7;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=7012;
 end   
19'd254714: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=39;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=8582;
 end   
19'd254715: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=3;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd254716: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=40;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd254717: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd254859: begin  
rid<=1;
end
19'd254860: begin  
end
19'd254861: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd254862: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd254863: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd254864: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd254865: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd254866: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd254867: begin  
rid<=0;
end
19'd255001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=80;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=17667;
 end   
19'd255002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=11;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11912;
 end   
19'd255003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=26;
   mapp<=50;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=15997;
 end   
19'd255004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=80;
   mapp<=66;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=14301;
 end   
19'd255005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=50;
   mapp<=95;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=17183;
 end   
19'd255006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=22;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd255007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=51;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd255008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=9;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd255009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=95;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd255010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=21;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=33510;
 end   
19'd255011: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=87;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=25462;
 end   
19'd255012: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=3;
   mapp<=87;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=30264;
 end   
19'd255013: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=50;
   mapp<=89;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=29811;
 end   
19'd255014: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=83;
   mapp<=31;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=31620;
 end   
19'd255015: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=10;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd255016: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=44;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd255017: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=69;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd255018: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=76;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd255019: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd255161: begin  
rid<=1;
end
19'd255162: begin  
end
19'd255163: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd255164: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd255165: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd255166: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd255167: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd255168: begin  
rid<=0;
end
19'd255301: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=65;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8313;
 end   
19'd255302: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=65;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd255303: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=24;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd255304: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=37;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd255305: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=4;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd255306: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=86;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd255307: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=26;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd255308: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=61;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd255309: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=79;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd255310: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=70;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=25439;
 end   
19'd255311: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=50;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd255312: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=18;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd255313: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=23;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd255314: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=3;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd255315: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=78;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd255316: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=47;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd255317: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=4;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd255318: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=91;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd255319: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd255461: begin  
rid<=1;
end
19'd255462: begin  
end
19'd255463: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd255464: begin  
rid<=0;
end
19'd255601: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=85;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=23441;
 end   
19'd255602: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=13;
   mapp<=30;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=27857;
 end   
19'd255603: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=70;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd255604: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=79;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd255605: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=52;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd255606: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=94;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd255607: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=63;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd255608: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=75;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd255609: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=8;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd255610: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=33;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd255611: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd255612: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=72;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=48929;
 end   
19'd255613: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=29;
   mapp<=65;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=51803;
 end   
19'd255614: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=32;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd255615: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=52;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd255616: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=34;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd255617: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=99;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd255618: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=61;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd255619: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=80;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd255620: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=57;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd255621: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=60;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd255622: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd255623: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd255765: begin  
rid<=1;
end
19'd255766: begin  
end
19'd255767: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd255768: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd255769: begin  
rid<=0;
end
19'd255901: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=13;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13726;
 end   
19'd255902: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=96;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd255903: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=50;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd255904: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=88;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=26024;
 end   
19'd255905: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=79;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd255906: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=42;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd255907: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd256049: begin  
rid<=1;
end
19'd256050: begin  
end
19'd256051: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd256052: begin  
rid<=0;
end
19'd256201: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=88;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6248;
 end   
19'd256202: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=81;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5761;
 end   
19'd256203: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=89;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6339;
 end   
19'd256204: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=73;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5213;
 end   
19'd256205: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=23;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1673;
 end   
19'd256206: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=46;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=3316;
 end   
19'd256207: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=39;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=2829;
 end   
19'd256208: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=80;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=5750;
 end   
19'd256209: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=68;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=4908;
 end   
19'd256210: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=98;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=7048;
 end   
19'd256211: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=7;
   mapp<=0;
   pp<=100;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[10]<=597;
 end   
19'd256212: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=16;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7768;
 end   
19'd256213: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=68;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=12221;
 end   
19'd256214: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=95;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15364;
 end   
19'd256215: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=98;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=14523;
 end   
19'd256216: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=50;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=6423;
 end   
19'd256217: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=69;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=9871;
 end   
19'd256218: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=41;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=6724;
 end   
19'd256219: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=59;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=11355;
 end   
19'd256220: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=92;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=13648;
 end   
19'd256221: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=85;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=15123;
 end   
19'd256222: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=53;
   mapp<=0;
   pp<=100;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[10]<=5632;
 end   
19'd256223: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd256365: begin  
rid<=1;
end
19'd256366: begin  
end
19'd256367: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd256368: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd256369: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd256370: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd256371: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd256372: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd256373: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd256374: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd256375: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd256376: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd256377: begin  
check0<=expctdoutput[10]-outcheck0;
end
19'd256378: begin  
rid<=0;
end
19'd256501: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=82;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6556;
 end   
19'd256502: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=66;
   mapp<=31;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6644;
 end   
19'd256503: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=62;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9526;
 end   
19'd256504: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=67;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=11596;
 end   
19'd256505: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=92;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=8970;
 end   
19'd256506: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=21;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=3818;
 end   
19'd256507: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd256508: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=46;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8948;
 end   
19'd256509: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=4;
   mapp<=69;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=10094;
 end   
19'd256510: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=69;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=12920;
 end   
19'd256511: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=55;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=14158;
 end   
19'd256512: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=8;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=9394;
 end   
19'd256513: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=14;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=4698;
 end   
19'd256514: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd256515: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd256657: begin  
rid<=1;
end
19'd256658: begin  
end
19'd256659: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd256660: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd256661: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd256662: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd256663: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd256664: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd256665: begin  
rid<=0;
end
19'd256801: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=16;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2708;
 end   
19'd256802: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=51;
   mapp<=28;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1376;
 end   
19'd256803: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=18;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4082;
 end   
19'd256804: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=74;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=2438;
 end   
19'd256805: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=24;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=832;
 end   
19'd256806: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=8;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=3646;
 end   
19'd256807: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=68;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=5738;
 end   
19'd256808: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd256809: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=42;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8630;
 end   
19'd256810: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=62;
   mapp<=84;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8500;
 end   
19'd256811: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=58;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=10424;
 end   
19'd256812: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=63;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=9300;
 end   
19'd256813: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=68;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=4742;
 end   
19'd256814: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=17;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=8266;
 end   
19'd256815: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=63;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=10864;
 end   
19'd256816: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd256817: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd256959: begin  
rid<=1;
end
19'd256960: begin  
end
19'd256961: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd256962: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd256963: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd256964: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd256965: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd256966: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd256967: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd256968: begin  
rid<=0;
end
19'd257101: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=22;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1166;
 end   
19'd257102: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=27;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1441;
 end   
19'd257103: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=14;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=762;
 end   
19'd257104: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=47;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=1213;
 end   
19'd257105: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=1;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=1442;
 end   
19'd257106: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=78;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=840;
 end   
19'd257107: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd257249: begin  
rid<=1;
end
19'd257250: begin  
end
19'd257251: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd257252: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd257253: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd257254: begin  
rid<=0;
end
19'd257401: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=78;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4760;
 end   
19'd257402: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=17;
   mapp<=18;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5062;
 end   
19'd257403: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=40;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd257404: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=22;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd257405: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=0;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd257406: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=93;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17021;
 end   
19'd257407: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=61;
   mapp<=18;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=13817;
 end   
19'd257408: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=67;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd257409: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=8;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd257410: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=0;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd257411: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd257553: begin  
rid<=1;
end
19'd257554: begin  
end
19'd257555: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd257556: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd257557: begin  
rid<=0;
end
19'd257701: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=60;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4200;
 end   
19'd257702: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=13;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=920;
 end   
19'd257703: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=78;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5480;
 end   
19'd257704: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=94;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6610;
 end   
19'd257705: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=86;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6060;
 end   
19'd257706: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=69;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=4880;
 end   
19'd257707: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=39;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=2790;
 end   
19'd257708: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=41;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=2940;
 end   
19'd257709: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=92;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=6520;
 end   
19'd257710: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=29;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=2120;
 end   
19'd257711: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=58;
   mapp<=0;
   pp<=100;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[10]<=4160;
 end   
19'd257712: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=82;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7398;
 end   
19'd257713: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=17;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=1583;
 end   
19'd257714: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=20;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=6260;
 end   
19'd257715: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=8;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6922;
 end   
19'd257716: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=42;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=7698;
 end   
19'd257717: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=14;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=5426;
 end   
19'd257718: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=4;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=2946;
 end   
19'd257719: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=35;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=4305;
 end   
19'd257720: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=39;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=8041;
 end   
19'd257721: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=4;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=2276;
 end   
19'd257722: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=65;
   mapp<=0;
   pp<=100;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[10]<=6695;
 end   
19'd257723: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd257865: begin  
rid<=1;
end
19'd257866: begin  
end
19'd257867: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd257868: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd257869: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd257870: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd257871: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd257872: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd257873: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd257874: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd257875: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd257876: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd257877: begin  
check0<=expctdoutput[10]-outcheck0;
end
19'd257878: begin  
rid<=0;
end
19'd258001: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=55;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16540;
 end   
19'd258002: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=83;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd258003: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=43;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd258004: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=86;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd258005: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=92;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd258006: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=82;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd258007: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=16;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd258008: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=34;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd258009: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=93;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd258010: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=27;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd258011: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=21;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=45189;
 end   
19'd258012: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=99;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd258013: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=40;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd258014: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=3;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd258015: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=98;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd258016: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=1;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd258017: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=86;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd258018: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=94;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd258019: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=61;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd258020: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=80;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd258021: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd258163: begin  
rid<=1;
end
19'd258164: begin  
end
19'd258165: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd258166: begin  
rid<=0;
end
19'd258301: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=62;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7189;
 end   
19'd258302: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=71;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6240;
 end   
19'd258303: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=61;
   mapp<=6;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2532;
 end   
19'd258304: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=17;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3242;
 end   
19'd258305: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=31;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6141;
 end   
19'd258306: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=64;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=5612;
 end   
19'd258307: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=54;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=3094;
 end   
19'd258308: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=20;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=8358;
 end   
19'd258309: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=94;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=4297;
 end   
19'd258310: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=31;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd258311: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=39;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd258312: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=92;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=18033;
 end   
19'd258313: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=44;
   mapp<=62;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=13578;
 end   
19'd258314: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=22;
   mapp<=26;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=10654;
 end   
19'd258315: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=91;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=13564;
 end   
19'd258316: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=26;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=12133;
 end   
19'd258317: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=48;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=11890;
 end   
19'd258318: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=34;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=8754;
 end   
19'd258319: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=9;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=16642;
 end   
19'd258320: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=89;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=17523;
 end   
19'd258321: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=78;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd258322: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=42;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd258323: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd258465: begin  
rid<=1;
end
19'd258466: begin  
end
19'd258467: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd258468: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd258469: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd258470: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd258471: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd258472: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd258473: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd258474: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd258475: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd258476: begin  
rid<=0;
end
19'd258601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=97;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=31747;
 end   
19'd258602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=32;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=26039;
 end   
19'd258603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=83;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd258604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=61;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd258605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=20;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd258606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=79;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd258607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=95;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd258608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=28;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd258609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd258610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=88;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=58903;
 end   
19'd258611: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=56;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=59369;
 end   
19'd258612: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=18;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd258613: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=84;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd258614: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=39;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd258615: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=74;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd258616: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=81;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd258617: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=64;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd258618: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd258619: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd258761: begin  
rid<=1;
end
19'd258762: begin  
end
19'd258763: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd258764: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd258765: begin  
rid<=0;
end
19'd258901: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=61;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14498;
 end   
19'd258902: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=45;
   mapp<=50;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=16721;
 end   
19'd258903: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=80;
   mapp<=45;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=16916;
 end   
19'd258904: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=41;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd258905: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=61;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd258906: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=7;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd258907: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=57;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd258908: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=43;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd258909: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=76;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd258910: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=92;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=33963;
 end   
19'd258911: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=52;
   mapp<=4;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=32612;
 end   
19'd258912: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=60;
   mapp<=63;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=31212;
 end   
19'd258913: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=77;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd258914: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=41;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd258915: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=22;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd258916: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=7;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd258917: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=73;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd258918: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=63;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd258919: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd259061: begin  
rid<=1;
end
19'd259062: begin  
end
19'd259063: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd259064: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd259065: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd259066: begin  
rid<=0;
end
19'd259201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=83;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=332;
 end   
19'd259202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=50;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4160;
 end   
19'd259203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=58;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4834;
 end   
19'd259204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=60;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5010;
 end   
19'd259205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=38;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=3866;
 end   
19'd259206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=53;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=6174;
 end   
19'd259207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=58;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=7038;
 end   
19'd259208: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=93;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=8544;
 end   
19'd259209: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd259351: begin  
rid<=1;
end
19'd259352: begin  
end
19'd259353: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd259354: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd259355: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd259356: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd259357: begin  
rid<=0;
end
19'd259501: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=16;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8471;
 end   
19'd259502: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=60;
   mapp<=12;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12427;
 end   
19'd259503: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=75;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd259504: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd259505: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=99;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17411;
 end   
19'd259506: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=21;
   mapp<=25;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=25252;
 end   
19'd259507: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=99;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd259508: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd259509: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd259651: begin  
rid<=1;
end
19'd259652: begin  
end
19'd259653: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd259654: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd259655: begin  
rid<=0;
end
19'd259801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=78;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7836;
 end   
19'd259802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=6;
   mapp<=58;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3486;
 end   
19'd259803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=50;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7140;
 end   
19'd259804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=40;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5552;
 end   
19'd259805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=29;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3868;
 end   
19'd259806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=18;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=2068;
 end   
19'd259807: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=5;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=2744;
 end   
19'd259808: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=38;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=7140;
 end   
19'd259809: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=59;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=8702;
 end   
19'd259810: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=51;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd259811: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=9;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=9678;
 end   
19'd259812: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=32;
   mapp<=30;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=9502;
 end   
19'd259813: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=96;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=18798;
 end   
19'd259814: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=75;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=14672;
 end   
19'd259815: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=59;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=11990;
 end   
19'd259816: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=78;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=11062;
 end   
19'd259817: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=45;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=8144;
 end   
19'd259818: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=33;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=12174;
 end   
19'd259819: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=60;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=15272;
 end   
19'd259820: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd259821: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd259963: begin  
rid<=1;
end
19'd259964: begin  
end
19'd259965: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd259966: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd259967: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd259968: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd259969: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd259970: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd259971: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd259972: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd259973: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd259974: begin  
rid<=0;
end
19'd260101: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=51;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4297;
 end   
19'd260102: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=47;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3769;
 end   
19'd260103: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=42;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6251;
 end   
19'd260104: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=87;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6864;
 end   
19'd260105: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=51;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5414;
 end   
19'd260106: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd260107: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=36;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8643;
 end   
19'd260108: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=49;
   mapp<=74;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=9765;
 end   
19'd260109: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=68;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=11149;
 end   
19'd260110: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=50;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=9154;
 end   
19'd260111: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=10;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=7146;
 end   
19'd260112: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd260113: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd260255: begin  
rid<=1;
end
19'd260256: begin  
end
19'd260257: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd260258: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd260259: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd260260: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd260261: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd260262: begin  
rid<=0;
end
19'd260401: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=10;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13649;
 end   
19'd260402: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=47;
   mapp<=13;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12358;
 end   
19'd260403: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=83;
   mapp<=32;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=18847;
 end   
19'd260404: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=46;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd260405: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=21;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd260406: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=57;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd260407: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=93;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd260408: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd260409: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd260410: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=22204;
 end   
19'd260411: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=97;
   mapp<=21;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=25308;
 end   
19'd260412: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=36;
   mapp<=50;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=36546;
 end   
19'd260413: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=36;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd260414: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=1;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd260415: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=11;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd260416: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=53;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd260417: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd260418: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd260419: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd260561: begin  
rid<=1;
end
19'd260562: begin  
end
19'd260563: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd260564: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd260565: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd260566: begin  
rid<=0;
end
19'd260701: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=95;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11491;
 end   
19'd260702: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=5;
   mapp<=78;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9643;
 end   
19'd260703: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=78;
   mapp<=72;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12872;
 end   
19'd260704: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=11;
   mapp<=15;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=9277;
 end   
19'd260705: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=63;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=9032;
 end   
19'd260706: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=93;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=14700;
 end   
19'd260707: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=23;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=5525;
 end   
19'd260708: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=68;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=7657;
 end   
19'd260709: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd260710: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd260711: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd260712: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=69;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=18205;
 end   
19'd260713: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=27;
   mapp<=21;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=14017;
 end   
19'd260714: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=47;
   mapp<=79;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=22442;
 end   
19'd260715: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=40;
   mapp<=16;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=17805;
 end   
19'd260716: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=1;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=16824;
 end   
19'd260717: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=91;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=28445;
 end   
19'd260718: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=78;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=17116;
 end   
19'd260719: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=40;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=17348;
 end   
19'd260720: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd260721: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd260722: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd260723: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd260865: begin  
rid<=1;
end
19'd260866: begin  
end
19'd260867: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd260868: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd260869: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd260870: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd260871: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd260872: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd260873: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd260874: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd260875: begin  
rid<=0;
end
19'd261001: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=5;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=921;
 end   
19'd261002: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=23;
   mapp<=27;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2238;
 end   
19'd261003: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=91;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1786;
 end   
19'd261004: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=57;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1603;
 end   
19'd261005: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=56;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=688;
 end   
19'd261006: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=16;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=1970;
 end   
19'd261007: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=80;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=966;
 end   
19'd261008: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=22;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=249;
 end   
19'd261009: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=3;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=877;
 end   
19'd261010: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd261011: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=22;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=1481;
 end   
19'd261012: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=15;
   mapp<=8;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=2444;
 end   
19'd261013: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=2;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=2280;
 end   
19'd261014: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=30;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=2743;
 end   
19'd261015: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=32;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=1422;
 end   
19'd261016: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=2;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=2704;
 end   
19'd261017: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=46;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=2248;
 end   
19'd261018: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=18;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=825;
 end   
19'd261019: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=12;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=2446;
 end   
19'd261020: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd261021: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd261163: begin  
rid<=1;
end
19'd261164: begin  
end
19'd261165: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd261166: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd261167: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd261168: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd261169: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd261170: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd261171: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd261172: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd261173: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd261174: begin  
rid<=0;
end
19'd261301: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=15;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13171;
 end   
19'd261302: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=65;
   mapp<=51;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=14913;
 end   
19'd261303: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=61;
   mapp<=99;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12359;
 end   
19'd261304: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=41;
   mapp<=92;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=10177;
 end   
19'd261305: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=51;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=8055;
 end   
19'd261306: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=43;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6038;
 end   
19'd261307: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=69;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=4267;
 end   
19'd261308: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=6;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=5753;
 end   
19'd261309: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd261310: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd261311: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd261312: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=23;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=29385;
 end   
19'd261313: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=87;
   mapp<=78;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=27159;
 end   
19'd261314: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=99;
   mapp<=72;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=26285;
 end   
19'd261315: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=91;
   mapp<=23;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=21807;
 end   
19'd261316: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=21;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=19585;
 end   
19'd261317: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=90;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=17986;
 end   
19'd261318: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=4;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=18817;
 end   
19'd261319: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=31;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=17973;
 end   
19'd261320: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd261321: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd261322: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd261323: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd261465: begin  
rid<=1;
end
19'd261466: begin  
end
19'd261467: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd261468: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd261469: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd261470: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd261471: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd261472: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd261473: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd261474: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd261475: begin  
rid<=0;
end
19'd261601: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=12;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=15442;
 end   
19'd261602: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=59;
   mapp<=52;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=14607;
 end   
19'd261603: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=97;
   mapp<=83;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8733;
 end   
19'd261604: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=49;
   mapp<=87;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=8429;
 end   
19'd261605: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=13;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=13174;
 end   
19'd261606: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=27;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=12333;
 end   
19'd261607: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=81;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=8118;
 end   
19'd261608: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd261609: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd261610: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd261611: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=68;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=28252;
 end   
19'd261612: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=41;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=22907;
 end   
19'd261613: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=87;
   mapp<=40;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=13751;
 end   
19'd261614: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=3;
   mapp<=3;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=9805;
 end   
19'd261615: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=25;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=19320;
 end   
19'd261616: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=19670;
 end   
19'd261617: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=49;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=14776;
 end   
19'd261618: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd261619: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd261620: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd261621: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd261763: begin  
rid<=1;
end
19'd261764: begin  
end
19'd261765: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd261766: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd261767: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd261768: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd261769: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd261770: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd261771: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd261772: begin  
rid<=0;
end
19'd261901: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=48;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3264;
 end   
19'd261902: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=53;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3614;
 end   
19'd261903: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=41;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=3346;
 end   
19'd261904: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=52;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=3718;
 end   
19'd261905: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd262047: begin  
rid<=1;
end
19'd262048: begin  
end
19'd262049: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd262050: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd262051: begin  
rid<=0;
end
19'd262201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=73;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9913;
 end   
19'd262202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=62;
   mapp<=41;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8605;
 end   
19'd262203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=85;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6109;
 end   
19'd262204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=57;
   mapp<=7;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3081;
 end   
19'd262205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=36;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5053;
 end   
19'd262206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=6;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=9169;
 end   
19'd262207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=51;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=5281;
 end   
19'd262208: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=99;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=5101;
 end   
19'd262209: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=2;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd262210: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=44;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd262211: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=69;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd262212: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=12;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12492;
 end   
19'd262213: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=64;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=11504;
 end   
19'd262214: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=12;
   mapp<=24;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=13307;
 end   
19'd262215: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=41;
   mapp<=31;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=11897;
 end   
19'd262216: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=37;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=16041;
 end   
19'd262217: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=86;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=22645;
 end   
19'd262218: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=29;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=14947;
 end   
19'd262219: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=53;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=18804;
 end   
19'd262220: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=98;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd262221: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=47;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd262222: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=58;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd262223: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd262365: begin  
rid<=1;
end
19'd262366: begin  
end
19'd262367: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd262368: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd262369: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd262370: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd262371: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd262372: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd262373: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd262374: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd262375: begin  
rid<=0;
end
19'd262501: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=89;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11098;
 end   
19'd262502: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=29;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd262503: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=96;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd262504: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=41;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd262505: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=6;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd262506: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=1;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd262507: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=49;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=23055;
 end   
19'd262508: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=47;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd262509: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=19;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd262510: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=4;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd262511: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=62;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd262512: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=63;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd262513: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd262655: begin  
rid<=1;
end
19'd262656: begin  
end
19'd262657: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd262658: begin  
rid<=0;
end
19'd262801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=68;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6048;
 end   
19'd262802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=99;
   mapp<=24;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7276;
 end   
19'd262803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=80;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6092;
 end   
19'd262804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=73;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5940;
 end   
19'd262805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=82;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd262806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=70;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=13646;
 end   
19'd262807: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=41;
   mapp<=88;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18149;
 end   
19'd262808: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=97;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=13469;
 end   
19'd262809: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=21;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=14705;
 end   
19'd262810: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=86;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd262811: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd262953: begin  
rid<=1;
end
19'd262954: begin  
end
19'd262955: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd262956: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd262957: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd262958: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd262959: begin  
rid<=0;
end
19'd263101: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=49;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1715;
 end   
19'd263102: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=41;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2019;
 end   
19'd263103: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=86;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4234;
 end   
19'd263104: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=80;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3950;
 end   
19'd263105: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=23;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1167;
 end   
19'd263106: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=43;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=2157;
 end   
19'd263107: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=17;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=1868;
 end   
19'd263108: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=2053;
 end   
19'd263109: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=73;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=5475;
 end   
19'd263110: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=59;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=4953;
 end   
19'd263111: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=17;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=1456;
 end   
19'd263112: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=83;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=3568;
 end   
19'd263113: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd263255: begin  
rid<=1;
end
19'd263256: begin  
end
19'd263257: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd263258: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd263259: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd263260: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd263261: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd263262: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd263263: begin  
rid<=0;
end
19'd263401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=14;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5833;
 end   
19'd263402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=30;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd263403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=63;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd263404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=93;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16447;
 end   
19'd263405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=82;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd263406: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=77;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd263407: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd263549: begin  
rid<=1;
end
19'd263550: begin  
end
19'd263551: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd263552: begin  
rid<=0;
end
19'd263701: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=15;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10586;
 end   
19'd263702: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=37;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11479;
 end   
19'd263703: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=86;
   mapp<=72;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11747;
 end   
19'd263704: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=6;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd263705: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=6;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd263706: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd263707: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=71;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd263708: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=6;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=19874;
 end   
19'd263709: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=90;
   mapp<=42;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=25062;
 end   
19'd263710: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=31;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=22842;
 end   
19'd263711: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=65;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd263712: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=55;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd263713: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=78;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd263714: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=81;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd263715: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd263857: begin  
rid<=1;
end
19'd263858: begin  
end
19'd263859: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd263860: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd263861: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd263862: begin  
rid<=0;
end
19'd264001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=30;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6010;
 end   
19'd264002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=44;
   mapp<=3;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7026;
 end   
19'd264003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=82;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd264004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=22;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd264005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=0;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd264006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=36;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=9178;
 end   
19'd264007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=14;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=13702;
 end   
19'd264008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=36;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd264009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=48;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd264010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=0;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd264011: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd264153: begin  
rid<=1;
end
19'd264154: begin  
end
19'd264155: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd264156: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd264157: begin  
rid<=0;
end
19'd264301: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=33;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7970;
 end   
19'd264302: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=7;
   mapp<=76;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10659;
 end   
19'd264303: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=48;
   mapp<=12;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=14471;
 end   
19'd264304: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=62;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd264305: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=71;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd264306: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=77;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd264307: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=42;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=15571;
 end   
19'd264308: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=52;
   mapp<=73;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20882;
 end   
19'd264309: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=83;
   mapp<=18;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=21820;
 end   
19'd264310: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=25;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd264311: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=54;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd264312: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=49;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd264313: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd264455: begin  
rid<=1;
end
19'd264456: begin  
end
19'd264457: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd264458: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd264459: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd264460: begin  
rid<=0;
end
19'd264601: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=89;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10719;
 end   
19'd264602: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=65;
   mapp<=3;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4066;
 end   
19'd264603: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=43;
   mapp<=26;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7384;
 end   
19'd264604: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=19;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd264605: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd264606: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd264607: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=62;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=22316;
 end   
19'd264608: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=87;
   mapp<=60;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18770;
 end   
19'd264609: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=43;
   mapp<=62;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=23939;
 end   
19'd264610: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=43;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd264611: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd264612: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd264613: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd264755: begin  
rid<=1;
end
19'd264756: begin  
end
19'd264757: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd264758: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd264759: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd264760: begin  
rid<=0;
end
19'd264901: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=60;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=15273;
 end   
19'd264902: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=34;
   mapp<=87;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=19566;
 end   
19'd264903: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=95;
   mapp<=31;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=19795;
 end   
19'd264904: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=24;
   mapp<=56;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=20559;
 end   
19'd264905: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=43;
   mapp<=90;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=20124;
 end   
19'd264906: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=17;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd264907: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=45;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd264908: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd264909: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd264910: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd264911: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd264912: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=80;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=40765;
 end   
19'd264913: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=3;
   mapp<=96;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=39862;
 end   
19'd264914: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=76;
   mapp<=96;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=38714;
 end   
19'd264915: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=52;
   mapp<=5;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=37825;
 end   
19'd264916: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=36;
   mapp<=38;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=40152;
 end   
19'd264917: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=98;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd264918: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=12;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd264919: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd264920: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd264921: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd264922: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd264923: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd265065: begin  
rid<=1;
end
19'd265066: begin  
end
19'd265067: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd265068: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd265069: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd265070: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd265071: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd265072: begin  
rid<=0;
end
19'd265201: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=23;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8914;
 end   
19'd265202: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=27;
   mapp<=89;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7703;
 end   
19'd265203: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=56;
   mapp<=73;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9461;
 end   
19'd265204: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=2;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd265205: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=20;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd265206: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd265207: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=65;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd265208: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=64;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=24119;
 end   
19'd265209: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=16;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=25459;
 end   
19'd265210: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=96;
   mapp<=75;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=24885;
 end   
19'd265211: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=77;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd265212: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=47;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd265213: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=19;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd265214: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=28;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd265215: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd265357: begin  
rid<=1;
end
19'd265358: begin  
end
19'd265359: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd265360: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd265361: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd265362: begin  
rid<=0;
end
19'd265501: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=33;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7898;
 end   
19'd265502: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=98;
   mapp<=21;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12993;
 end   
19'd265503: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=59;
   mapp<=14;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12998;
 end   
19'd265504: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=78;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd265505: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=19;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd265506: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=79;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd265507: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=84;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd265508: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=93;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=28309;
 end   
19'd265509: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=86;
   mapp<=28;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=25634;
 end   
19'd265510: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=78;
   mapp<=93;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=26380;
 end   
19'd265511: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=43;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd265512: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=80;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd265513: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=6;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd265514: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd265515: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd265657: begin  
rid<=1;
end
19'd265658: begin  
end
19'd265659: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd265660: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd265661: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd265662: begin  
rid<=0;
end
19'd265801: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=18;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4319;
 end   
19'd265802: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=17;
   mapp<=99;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4212;
 end   
19'd265803: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=14;
   mapp<=88;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3706;
 end   
19'd265804: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=66;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3276;
 end   
19'd265805: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=70;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2494;
 end   
19'd265806: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=62;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=1462;
 end   
19'd265807: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=10;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=1065;
 end   
19'd265808: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=9;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=2392;
 end   
19'd265809: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=48;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=3556;
 end   
19'd265810: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd265811: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd265812: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=99;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=11705;
 end   
19'd265813: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=78;
   mapp<=37;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=13935;
 end   
19'd265814: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=18;
   mapp<=74;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=13828;
 end   
19'd265815: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=16;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=12126;
 end   
19'd265816: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=86;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=14650;
 end   
19'd265817: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=31;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=10699;
 end   
19'd265818: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=68;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=12369;
 end   
19'd265819: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=48;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=11740;
 end   
19'd265820: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=46;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=13612;
 end   
19'd265821: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd265822: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd265823: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd265965: begin  
rid<=1;
end
19'd265966: begin  
end
19'd265967: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd265968: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd265969: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd265970: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd265971: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd265972: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd265973: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd265974: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd265975: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd265976: begin  
rid<=0;
end
19'd266101: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=27;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9751;
 end   
19'd266102: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=88;
   mapp<=98;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6732;
 end   
19'd266103: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=13;
   mapp<=41;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5569;
 end   
19'd266104: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=36;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=10705;
 end   
19'd266105: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=98;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=10172;
 end   
19'd266106: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=83;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=4537;
 end   
19'd266107: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=14;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=8043;
 end   
19'd266108: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=78;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=7881;
 end   
19'd266109: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd266110: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd266111: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=14;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=10387;
 end   
19'd266112: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=14;
   mapp<=3;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=7359;
 end   
19'd266113: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=3;
   mapp<=30;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=6774;
 end   
19'd266114: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=55;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=11668;
 end   
19'd266115: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=5;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=11047;
 end   
19'd266116: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=41;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=6324;
 end   
19'd266117: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=77;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=10015;
 end   
19'd266118: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=45;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=9872;
 end   
19'd266119: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd266120: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd266121: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd266263: begin  
rid<=1;
end
19'd266264: begin  
end
19'd266265: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd266266: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd266267: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd266268: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd266269: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd266270: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd266271: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd266272: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd266273: begin  
rid<=0;
end
19'd266401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=63;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9630;
 end   
19'd266402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=90;
   mapp<=29;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5295;
 end   
19'd266403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=90;
   mapp<=71;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5550;
 end   
19'd266404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=25;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5496;
 end   
19'd266405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=55;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2495;
 end   
19'd266406: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=51;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=4071;
 end   
19'd266407: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=6;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd266408: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=47;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd266409: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=39;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17864;
 end   
19'd266410: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=28;
   mapp<=22;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=9439;
 end   
19'd266411: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=59;
   mapp<=65;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15152;
 end   
19'd266412: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=2;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=12643;
 end   
19'd266413: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=59;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=14942;
 end   
19'd266414: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=87;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=14333;
 end   
19'd266415: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=74;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd266416: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=3;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd266417: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd266559: begin  
rid<=1;
end
19'd266560: begin  
end
19'd266561: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd266562: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd266563: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd266564: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd266565: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd266566: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd266567: begin  
rid<=0;
end
19'd266701: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=57;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11639;
 end   
19'd266702: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=25;
   mapp<=31;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11822;
 end   
19'd266703: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=16;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd266704: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=79;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd266705: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=12;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd266706: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=95;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd266707: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd266708: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=79;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17683;
 end   
19'd266709: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=48;
   mapp<=7;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20274;
 end   
19'd266710: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=4;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd266711: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=20;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd266712: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=53;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd266713: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=41;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd266714: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd266715: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd266857: begin  
rid<=1;
end
19'd266858: begin  
end
19'd266859: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd266860: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd266861: begin  
rid<=0;
end
19'd267001: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=51;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1141;
 end   
19'd267002: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=86;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd267003: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=55;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=4702;
 end   
19'd267004: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=48;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd267005: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd267147: begin  
rid<=1;
end
19'd267148: begin  
end
19'd267149: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd267150: begin  
rid<=0;
end
19'd267301: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=91;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5999;
 end   
19'd267302: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=61;
   mapp<=70;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1519;
 end   
19'd267303: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=5;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=465;
 end   
19'd267304: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=5;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3555;
 end   
19'd267305: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=49;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4261;
 end   
19'd267306: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=47;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=5493;
 end   
19'd267307: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=65;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=6895;
 end   
19'd267308: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=80;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd267309: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=93;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=6464;
 end   
19'd267310: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=0;
   mapp<=61;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=3837;
 end   
19'd267311: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=38;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=2241;
 end   
19'd267312: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=26;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=7772;
 end   
19'd267313: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=67;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=9781;
 end   
19'd267314: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=85;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=7504;
 end   
19'd267315: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=26;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=12393;
 end   
19'd267316: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd267317: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd267459: begin  
rid<=1;
end
19'd267460: begin  
end
19'd267461: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd267462: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd267463: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd267464: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd267465: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd267466: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd267467: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd267468: begin  
rid<=0;
end
19'd267601: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=99;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13286;
 end   
19'd267602: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=78;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd267603: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=83;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd267604: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=60;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd267605: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=70;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16336;
 end   
19'd267606: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=13;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd267607: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=18;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd267608: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=4;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd267609: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd267751: begin  
rid<=1;
end
19'd267752: begin  
end
19'd267753: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd267754: begin  
rid<=0;
end
19'd267901: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=26;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=988;
 end   
19'd267902: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=71;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2708;
 end   
19'd267903: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=84;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3212;
 end   
19'd267904: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=42;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1626;
 end   
19'd267905: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=92;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3536;
 end   
19'd267906: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=53;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5228;
 end   
19'd267907: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=3;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=2948;
 end   
19'd267908: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=25;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=5212;
 end   
19'd267909: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=96;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=9306;
 end   
19'd267910: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=80;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=9936;
 end   
19'd267911: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd268053: begin  
rid<=1;
end
19'd268054: begin  
end
19'd268055: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd268056: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd268057: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd268058: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd268059: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd268060: begin  
rid<=0;
end
19'd268201: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=94;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1692;
 end   
19'd268202: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=480;
 end   
19'd268203: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=23;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2182;
 end   
19'd268204: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=75;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7080;
 end   
19'd268205: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=49;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4646;
 end   
19'd268206: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=82;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7758;
 end   
19'd268207: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=60;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=5700;
 end   
19'd268208: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=96;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5436;
 end   
19'd268209: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=65;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=6720;
 end   
19'd268210: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=93;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=11110;
 end   
19'd268211: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=57;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=12552;
 end   
19'd268212: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=68;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=11174;
 end   
19'd268213: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=34;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=11022;
 end   
19'd268214: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=29;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=8484;
 end   
19'd268215: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd268357: begin  
rid<=1;
end
19'd268358: begin  
end
19'd268359: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd268360: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd268361: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd268362: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd268363: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd268364: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd268365: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd268366: begin  
rid<=0;
end
19'd268501: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=57;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9498;
 end   
19'd268502: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=33;
   mapp<=33;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11305;
 end   
19'd268503: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=33;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=14675;
 end   
19'd268504: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=9;
   mapp<=1;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=11085;
 end   
19'd268505: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=93;
   mapp<=52;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=13342;
 end   
19'd268506: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd268507: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd268508: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd268509: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd268510: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=17;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17420;
 end   
19'd268511: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=34;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=17655;
 end   
19'd268512: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=99;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=19376;
 end   
19'd268513: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=19;
   mapp<=3;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=17388;
 end   
19'd268514: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=92;
   mapp<=0;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=18287;
 end   
19'd268515: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd268516: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd268517: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd268518: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd268519: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd268661: begin  
rid<=1;
end
19'd268662: begin  
end
19'd268663: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd268664: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd268665: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd268666: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd268667: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd268668: begin  
rid<=0;
end
19'd268801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=49;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4704;
 end   
19'd268802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=0;
   mapp<=85;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4175;
 end   
19'd268803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=77;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=10787;
 end   
19'd268804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=0;
   mapp<=36;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=6947;
 end   
19'd268805: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd268947: begin  
rid<=1;
end
19'd268948: begin  
end
19'd268949: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd268950: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd268951: begin  
rid<=0;
end
19'd269101: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=16;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=23546;
 end   
19'd269102: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=60;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd269103: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=94;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd269104: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=88;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd269105: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=42;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd269106: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=73;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd269107: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=20;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd269108: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=22;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd269109: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=60;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd269110: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=56;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd269111: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=21;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=36572;
 end   
19'd269112: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=95;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd269113: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=55;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd269114: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=40;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd269115: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=11;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd269116: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=18;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd269117: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=23;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd269118: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=7;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd269119: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=39;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd269120: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=39;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd269121: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd269263: begin  
rid<=1;
end
19'd269264: begin  
end
19'd269265: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd269266: begin  
rid<=0;
end
19'd269401: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=95;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10122;
 end   
19'd269402: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=53;
   mapp<=44;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7211;
 end   
19'd269403: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=57;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5594;
 end   
19'd269404: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=3;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1746;
 end   
19'd269405: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=27;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=7110;
 end   
19'd269406: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=85;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=10616;
 end   
19'd269407: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=47;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=6062;
 end   
19'd269408: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=29;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=5157;
 end   
19'd269409: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=44;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=6274;
 end   
19'd269410: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd269411: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=97;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=18719;
 end   
19'd269412: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=69;
   mapp<=29;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=14923;
 end   
19'd269413: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=71;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=15310;
 end   
19'd269414: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=41;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=8690;
 end   
19'd269415: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=43;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=13834;
 end   
19'd269416: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=37;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=20001;
 end   
19'd269417: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=84;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=14555;
 end   
19'd269418: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=5;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=10541;
 end   
19'd269419: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=71;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=13644;
 end   
19'd269420: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd269421: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd269563: begin  
rid<=1;
end
19'd269564: begin  
end
19'd269565: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd269566: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd269567: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd269568: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd269569: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd269570: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd269571: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd269572: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd269573: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd269574: begin  
rid<=0;
end
19'd269701: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=79;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14362;
 end   
19'd269702: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=70;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd269703: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=38;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd269704: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=68;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd269705: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=29;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd269706: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=56;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd269707: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=80;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=26959;
 end   
19'd269708: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=49;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd269709: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=25;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd269710: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=25;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd269711: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=4;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd269712: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=45;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd269713: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd269855: begin  
rid<=1;
end
19'd269856: begin  
end
19'd269857: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd269858: begin  
rid<=0;
end
19'd270001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=64;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13344;
 end   
19'd270002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=51;
   mapp<=39;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=14946;
 end   
19'd270003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=70;
   mapp<=69;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=13637;
 end   
19'd270004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=69;
   mapp<=89;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=15816;
 end   
19'd270005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=39;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=12678;
 end   
19'd270006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=28;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=11730;
 end   
19'd270007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=89;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=14602;
 end   
19'd270008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=36;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=9838;
 end   
19'd270009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd270010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd270011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd270012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=81;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=29634;
 end   
19'd270013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=51;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=30424;
 end   
19'd270014: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=33;
   mapp<=18;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=22910;
 end   
19'd270015: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=82;
   mapp<=78;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=27724;
 end   
19'd270016: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=79;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=23059;
 end   
19'd270017: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=15;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=21700;
 end   
19'd270018: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=13;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=27246;
 end   
19'd270019: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=34;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=22553;
 end   
19'd270020: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd270021: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd270022: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd270023: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd270165: begin  
rid<=1;
end
19'd270166: begin  
end
19'd270167: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd270168: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd270169: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd270170: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd270171: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd270172: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd270173: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd270174: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd270175: begin  
rid<=0;
end
19'd270301: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=28;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=22442;
 end   
19'd270302: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=71;
   mapp<=89;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15614;
 end   
19'd270303: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=88;
   mapp<=40;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=20874;
 end   
19'd270304: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=37;
   mapp<=60;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=12486;
 end   
19'd270305: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=15;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd270306: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=6;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd270307: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=99;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd270308: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=13;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd270309: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd270310: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd270311: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd270312: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=78;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=38488;
 end   
19'd270313: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=36;
   mapp<=23;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=30342;
 end   
19'd270314: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=5;
   mapp<=31;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=38058;
 end   
19'd270315: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=19;
   mapp<=55;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=25857;
 end   
19'd270316: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=10;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd270317: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=35;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd270318: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=60;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd270319: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=93;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd270320: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd270321: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd270322: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd270323: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd270465: begin  
rid<=1;
end
19'd270466: begin  
end
19'd270467: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd270468: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd270469: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd270470: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd270471: begin  
rid<=0;
end
19'd270601: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=23;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1587;
 end   
19'd270602: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=43;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=999;
 end   
19'd270603: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=23;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=549;
 end   
19'd270604: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=41;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=973;
 end   
19'd270605: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=1;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=63;
 end   
19'd270606: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=20;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=510;
 end   
19'd270607: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=84;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=1992;
 end   
19'd270608: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=70;
 end   
19'd270609: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=89;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=2127;
 end   
19'd270610: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=63;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=1539;
 end   
19'd270611: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=85;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=2862;
 end   
19'd270612: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=60;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=6099;
 end   
19'd270613: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=92;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=8369;
 end   
19'd270614: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=92;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=8793;
 end   
19'd270615: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=50;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=4313;
 end   
19'd270616: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=14;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=1700;
 end   
19'd270617: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=67;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=7687;
 end   
19'd270618: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=58;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=5000;
 end   
19'd270619: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=15;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=3402;
 end   
19'd270620: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=53;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=6044;
 end   
19'd270621: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd270763: begin  
rid<=1;
end
19'd270764: begin  
end
19'd270765: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd270766: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd270767: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd270768: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd270769: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd270770: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd270771: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd270772: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd270773: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd270774: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd270775: begin  
rid<=0;
end
19'd270901: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=80;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14476;
 end   
19'd270902: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=16;
   mapp<=59;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8240;
 end   
19'd270903: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=72;
   mapp<=86;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11872;
 end   
19'd270904: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=10;
   mapp<=22;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7552;
 end   
19'd270905: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=55;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6672;
 end   
19'd270906: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=66;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=8126;
 end   
19'd270907: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd270908: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd270909: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd270910: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd270911: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=79;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=19409;
 end   
19'd270912: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=4;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=13341;
 end   
19'd270913: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=42;
   mapp<=38;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=18892;
 end   
19'd270914: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=99;
   mapp<=12;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=16303;
 end   
19'd270915: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=37;
   mapp<=41;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=23266;
 end   
19'd270916: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=6;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=24662;
 end   
19'd270917: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd270918: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd270919: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd270920: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd270921: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd271063: begin  
rid<=1;
end
19'd271064: begin  
end
19'd271065: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd271066: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd271067: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd271068: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd271069: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd271070: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd271071: begin  
rid<=0;
end
19'd271201: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=57;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14767;
 end   
19'd271202: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=89;
   mapp<=71;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=14009;
 end   
19'd271203: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=49;
   mapp<=78;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=10991;
 end   
19'd271204: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=21;
   mapp<=52;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=8900;
 end   
19'd271205: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd271206: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd271207: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd271208: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=60;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=22043;
 end   
19'd271209: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=10;
   mapp<=1;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20427;
 end   
19'd271210: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=1;
   mapp<=50;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=19734;
 end   
19'd271211: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=64;
   mapp<=34;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=15261;
 end   
19'd271212: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd271213: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd271214: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd271215: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd271357: begin  
rid<=1;
end
19'd271358: begin  
end
19'd271359: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd271360: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd271361: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd271362: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd271363: begin  
rid<=0;
end
19'd271501: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=18;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=20152;
 end   
19'd271502: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=52;
   mapp<=21;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=19949;
 end   
19'd271503: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=40;
   mapp<=19;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=18886;
 end   
19'd271504: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=41;
   mapp<=86;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=17995;
 end   
19'd271505: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=66;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd271506: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=67;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd271507: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=64;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd271508: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=15;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd271509: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd271510: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd271511: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd271512: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=87;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=39415;
 end   
19'd271513: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=21;
   mapp<=42;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=35780;
 end   
19'd271514: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=38;
   mapp<=84;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=38002;
 end   
19'd271515: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=3;
   mapp<=18;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=25114;
 end   
19'd271516: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=67;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd271517: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=84;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd271518: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=95;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd271519: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=11;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd271520: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd271521: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd271522: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd271523: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd271665: begin  
rid<=1;
end
19'd271666: begin  
end
19'd271667: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd271668: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd271669: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd271670: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd271671: begin  
rid<=0;
end
19'd271801: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=12;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=420;
 end   
19'd271802: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=63;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=3759;
 end   
19'd271803: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd271945: begin  
rid<=1;
end
19'd271946: begin  
end
19'd271947: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd271948: begin  
rid<=0;
end
19'd272101: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=66;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14877;
 end   
19'd272102: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=48;
   mapp<=8;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11200;
 end   
19'd272103: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=14;
   mapp<=52;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=15009;
 end   
19'd272104: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=52;
   mapp<=27;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=19288;
 end   
19'd272105: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=32;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd272106: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=39;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd272107: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=81;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd272108: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=94;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd272109: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd272110: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd272111: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd272112: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=54;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=31913;
 end   
19'd272113: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=66;
   mapp<=31;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=37981;
 end   
19'd272114: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=28;
   mapp<=95;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=45597;
 end   
19'd272115: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=75;
   mapp<=32;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=47436;
 end   
19'd272116: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=86;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd272117: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd272118: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=10;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd272119: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=94;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd272120: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd272121: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd272122: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd272123: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd272265: begin  
rid<=1;
end
19'd272266: begin  
end
19'd272267: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd272268: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd272269: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd272270: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd272271: begin  
rid<=0;
end
19'd272401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=51;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16140;
 end   
19'd272402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=32;
   mapp<=61;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=18025;
 end   
19'd272403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=81;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd272404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=75;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd272405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=36;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd272406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=40;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd272407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=36;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd272408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=58;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd272409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=27;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd272410: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=2;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=31634;
 end   
19'd272411: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=91;
   mapp<=6;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=41875;
 end   
19'd272412: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=78;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd272413: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=27;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd272414: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=65;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd272415: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=48;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd272416: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=59;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd272417: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=88;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd272418: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=54;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd272419: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd272561: begin  
rid<=1;
end
19'd272562: begin  
end
19'd272563: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd272564: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd272565: begin  
rid<=0;
end
19'd272701: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=97;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=18333;
 end   
19'd272702: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=90;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15989;
 end   
19'd272703: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=73;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8541;
 end   
19'd272704: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=16;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=9412;
 end   
19'd272705: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd272706: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=38;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=21019;
 end   
19'd272707: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=71;
   mapp<=10;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=23043;
 end   
19'd272708: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=94;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=14882;
 end   
19'd272709: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=39;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=13166;
 end   
19'd272710: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd272711: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd272853: begin  
rid<=1;
end
19'd272854: begin  
end
19'd272855: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd272856: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd272857: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd272858: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd272859: begin  
rid<=0;
end
19'd273001: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=61;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8087;
 end   
19'd273002: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=26;
   mapp<=89;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9593;
 end   
19'd273003: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=62;
   mapp<=34;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6204;
 end   
19'd273004: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=59;
   mapp<=28;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6280;
 end   
19'd273005: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=26;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=9529;
 end   
19'd273006: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=30;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=13462;
 end   
19'd273007: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd273008: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd273009: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd273010: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=61;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12434;
 end   
19'd273011: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=15;
   mapp<=53;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=17710;
 end   
19'd273012: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=49;
   mapp<=9;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=12182;
 end   
19'd273013: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=22;
   mapp<=61;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=13382;
 end   
19'd273014: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=80;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=18287;
 end   
19'd273015: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=27;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=19217;
 end   
19'd273016: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd273017: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd273018: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd273019: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd273161: begin  
rid<=1;
end
19'd273162: begin  
end
19'd273163: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd273164: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd273165: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd273166: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd273167: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd273168: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd273169: begin  
rid<=0;
end
19'd273301: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=48;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10914;
 end   
19'd273302: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=42;
   mapp<=84;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=16255;
 end   
19'd273303: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=24;
   mapp<=98;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11036;
 end   
19'd273304: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=81;
   mapp<=10;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=9609;
 end   
19'd273305: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=97;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=14929;
 end   
19'd273306: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd273307: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd273308: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd273309: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=6;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=19102;
 end   
19'd273310: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=10;
   mapp<=63;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=25003;
 end   
19'd273311: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=70;
   mapp<=19;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=21997;
 end   
19'd273312: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=89;
   mapp<=66;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=23157;
 end   
19'd273313: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=40;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=30181;
 end   
19'd273314: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd273315: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd273316: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd273317: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd273459: begin  
rid<=1;
end
19'd273460: begin  
end
19'd273461: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd273462: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd273463: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd273464: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd273465: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd273466: begin  
rid<=0;
end
19'd273601: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=24;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=22789;
 end   
19'd273602: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=43;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd273603: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=82;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd273604: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=59;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd273605: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=35;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd273606: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=95;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd273607: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=51;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd273608: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=91;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd273609: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=42;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd273610: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=70;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd273611: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=62;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=51344;
 end   
19'd273612: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=26;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd273613: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=3;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd273614: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=59;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd273615: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=65;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd273616: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=87;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd273617: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=9;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd273618: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=88;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd273619: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=83;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd273620: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=91;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd273621: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd273763: begin  
rid<=1;
end
19'd273764: begin  
end
19'd273765: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd273766: begin  
rid<=0;
end
19'd273901: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=4;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9003;
 end   
19'd273902: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=41;
   mapp<=42;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5599;
 end   
19'd273903: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=85;
   mapp<=85;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5069;
 end   
19'd273904: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=17;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=10152;
 end   
19'd273905: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=37;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=8329;
 end   
19'd273906: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=98;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=10708;
 end   
19'd273907: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=43;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=10903;
 end   
19'd273908: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=88;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=6491;
 end   
19'd273909: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=77;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=3994;
 end   
19'd273910: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd273911: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=22;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd273912: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=90;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17083;
 end   
19'd273913: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=5;
   mapp<=28;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8409;
 end   
19'd273914: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=70;
   mapp<=80;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=12661;
 end   
19'd273915: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=9;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=18158;
 end   
19'd273916: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=69;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=16407;
 end   
19'd273917: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=73;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=15610;
 end   
19'd273918: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=53;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=18813;
 end   
19'd273919: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=19;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=15965;
 end   
19'd273920: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=75;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=8912;
 end   
19'd273921: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=86;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd273922: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=7;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd273923: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd274065: begin  
rid<=1;
end
19'd274066: begin  
end
19'd274067: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd274068: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd274069: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd274070: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd274071: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd274072: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd274073: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd274074: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd274075: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd274076: begin  
rid<=0;
end
19'd274201: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=65;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14089;
 end   
19'd274202: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=51;
   mapp<=42;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=13320;
 end   
19'd274203: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=36;
   mapp<=3;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11778;
 end   
19'd274204: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=54;
   mapp<=24;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=12179;
 end   
19'd274205: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=35;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd274206: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=76;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd274207: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=38;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd274208: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=81;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd274209: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd274210: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd274211: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd274212: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=50;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=32112;
 end   
19'd274213: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=36;
   mapp<=24;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=30246;
 end   
19'd274214: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=45;
   mapp<=32;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=29357;
 end   
19'd274215: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=21;
   mapp<=52;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=32054;
 end   
19'd274216: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=63;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd274217: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=94;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd274218: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=81;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd274219: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=39;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd274220: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd274221: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd274222: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd274223: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd274365: begin  
rid<=1;
end
19'd274366: begin  
end
19'd274367: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd274368: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd274369: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd274370: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd274371: begin  
rid<=0;
end
19'd274501: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=60;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5340;
 end   
19'd274502: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10;
 end   
19'd274503: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=77;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6873;
 end   
19'd274504: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=74;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6616;
 end   
19'd274505: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=33;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2977;
 end   
19'd274506: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=86;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7704;
 end   
19'd274507: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=55;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=4955;
 end   
19'd274508: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=79;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=7101;
 end   
19'd274509: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=13;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=6211;
 end   
19'd274510: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=55;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=3695;
 end   
19'd274511: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=89;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=12836;
 end   
19'd274512: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=95;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=12981;
 end   
19'd274513: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=43;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=5858;
 end   
19'd274514: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=12;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=8508;
 end   
19'd274515: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=4;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=5223;
 end   
19'd274516: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=79;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=12394;
 end   
19'd274517: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd274659: begin  
rid<=1;
end
19'd274660: begin  
end
19'd274661: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd274662: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd274663: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd274664: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd274665: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd274666: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd274667: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd274668: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd274669: begin  
rid<=0;
end
19'd274801: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=74;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=15353;
 end   
19'd274802: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=5;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd274803: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=48;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd274804: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=88;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd274805: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=77;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd274806: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=43;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=22174;
 end   
19'd274807: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=20;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd274808: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd274809: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=16;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd274810: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=82;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd274811: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd274953: begin  
rid<=1;
end
19'd274954: begin  
end
19'd274955: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd274956: begin  
rid<=0;
end
19'd275101: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=15;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=900;
 end   
19'd275102: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=75;
   mapp<=8;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3655;
 end   
19'd275103: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=47;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7700;
 end   
19'd275104: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=93;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3075;
 end   
19'd275105: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=22;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3970;
 end   
19'd275106: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=48;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=3245;
 end   
19'd275107: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=33;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=4455;
 end   
19'd275108: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=52;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=7450;
 end   
19'd275109: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=88;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=5225;
 end   
19'd275110: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd275111: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=5;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=2396;
 end   
19'd275112: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=16;
   mapp<=91;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=5278;
 end   
19'd275113: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=73;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=8289;
 end   
19'd275114: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=14;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=4329;
 end   
19'd275115: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=74;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=4420;
 end   
19'd275116: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=5;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=4662;
 end   
19'd275117: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=87;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=6266;
 end   
19'd275118: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=86;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=9368;
 end   
19'd275119: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=93;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=5882;
 end   
19'd275120: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd275121: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd275263: begin  
rid<=1;
end
19'd275264: begin  
end
19'd275265: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd275266: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd275267: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd275268: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd275269: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd275270: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd275271: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd275272: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd275273: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd275274: begin  
rid<=0;
end
19'd275401: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=53;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4293;
 end   
19'd275402: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=96;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7786;
 end   
19'd275403: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=87;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7067;
 end   
19'd275404: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=61;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4971;
 end   
19'd275405: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=14;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1174;
 end   
19'd275406: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=49;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=4019;
 end   
19'd275407: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=75;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=6135;
 end   
19'd275408: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=84;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8157;
 end   
19'd275409: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=48;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=9994;
 end   
19'd275410: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=33;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=8585;
 end   
19'd275411: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=17;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=5753;
 end   
19'd275412: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=78;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=4762;
 end   
19'd275413: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=12;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=4571;
 end   
19'd275414: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=34;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=7699;
 end   
19'd275415: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd275557: begin  
rid<=1;
end
19'd275558: begin  
end
19'd275559: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd275560: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd275561: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd275562: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd275563: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd275564: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd275565: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd275566: begin  
rid<=0;
end
19'd275701: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=58;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14116;
 end   
19'd275702: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=54;
   mapp<=66;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=14938;
 end   
19'd275703: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=77;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=17225;
 end   
19'd275704: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=72;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=18298;
 end   
19'd275705: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=80;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=15604;
 end   
19'd275706: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=94;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=10738;
 end   
19'd275707: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=32;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=4786;
 end   
19'd275708: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=3;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd275709: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=24;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd275710: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=20;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=21421;
 end   
19'd275711: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=93;
   mapp<=51;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=26653;
 end   
19'd275712: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=54;
   mapp<=13;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=24667;
 end   
19'd275713: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=24;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=26340;
 end   
19'd275714: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=92;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=29365;
 end   
19'd275715: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=86;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=22716;
 end   
19'd275716: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=63;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=13745;
 end   
19'd275717: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=59;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd275718: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=7;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd275719: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd275861: begin  
rid<=1;
end
19'd275862: begin  
end
19'd275863: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd275864: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd275865: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd275866: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd275867: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd275868: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd275869: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd275870: begin  
rid<=0;
end
19'd276001: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=93;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9769;
 end   
19'd276002: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=82;
   mapp<=25;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7866;
 end   
19'd276003: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=42;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5081;
 end   
19'd276004: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=63;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6784;
 end   
19'd276005: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=61;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=7203;
 end   
19'd276006: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=84;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=8672;
 end   
19'd276007: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=66;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=5938;
 end   
19'd276008: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=16;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=3823;
 end   
19'd276009: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=97;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=9756;
 end   
19'd276010: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=65;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd276011: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=51;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16117;
 end   
19'd276012: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=25;
   mapp<=54;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=13070;
 end   
19'd276013: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=51;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=11159;
 end   
19'd276014: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=20;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=13604;
 end   
19'd276015: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=90;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=18237;
 end   
19'd276016: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=41;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=17928;
 end   
19'd276017: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=97;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=17874;
 end   
19'd276018: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=45;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=10015;
 end   
19'd276019: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=33;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=13260;
 end   
19'd276020: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=5;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd276021: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd276163: begin  
rid<=1;
end
19'd276164: begin  
end
19'd276165: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd276166: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd276167: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd276168: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd276169: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd276170: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd276171: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd276172: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd276173: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd276174: begin  
rid<=0;
end
19'd276301: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=80;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1792;
 end   
19'd276302: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=27;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2141;
 end   
19'd276303: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=18;
   mapp<=21;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=4688;
 end   
19'd276304: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=78;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=8187;
 end   
19'd276305: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=49;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4977;
 end   
19'd276306: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=33;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=3347;
 end   
19'd276307: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=7;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=2978;
 end   
19'd276308: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd276309: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd276310: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=7;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=12881;
 end   
19'd276311: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=93;
   mapp<=69;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=10263;
 end   
19'd276312: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=86;
   mapp<=47;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=16377;
 end   
19'd276313: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=38;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=22162;
 end   
19'd276314: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=91;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=18339;
 end   
19'd276315: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=61;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=18538;
 end   
19'd276316: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=82;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=19183;
 end   
19'd276317: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd276318: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd276319: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd276461: begin  
rid<=1;
end
19'd276462: begin  
end
19'd276463: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd276464: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd276465: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd276466: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd276467: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd276468: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd276469: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd276470: begin  
rid<=0;
end
19'd276601: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=90;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4752;
 end   
19'd276602: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=33;
   mapp<=24;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2134;
 end   
19'd276603: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=28;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2524;
 end   
19'd276604: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=53;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4738;
 end   
19'd276605: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=99;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5452;
 end   
19'd276606: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=44;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=4290;
 end   
19'd276607: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=96;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=4284;
 end   
19'd276608: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=238;
 end   
19'd276609: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=7;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=676;
 end   
19'd276610: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=12;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=2466;
 end   
19'd276611: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=77;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd276612: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=32;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=7805;
 end   
19'd276613: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=15;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=5664;
 end   
19'd276614: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=67;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=9952;
 end   
19'd276615: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=61;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=10257;
 end   
19'd276616: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=20;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=7172;
 end   
19'd276617: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=4;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=6811;
 end   
19'd276618: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=63;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=10206;
 end   
19'd276619: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=27;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=5171;
 end   
19'd276620: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=80;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=8081;
 end   
19'd276621: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=31;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=8310;
 end   
19'd276622: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=97;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd276623: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd276765: begin  
rid<=1;
end
19'd276766: begin  
end
19'd276767: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd276768: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd276769: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd276770: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd276771: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd276772: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd276773: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd276774: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd276775: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd276776: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd276777: begin  
rid<=0;
end
19'd276901: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=70;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6284;
 end   
19'd276902: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=62;
   mapp<=37;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6911;
 end   
19'd276903: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=91;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7612;
 end   
19'd276904: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=65;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7324;
 end   
19'd276905: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=97;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=7234;
 end   
19'd276906: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=45;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=5908;
 end   
19'd276907: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd276908: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=70;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14164;
 end   
19'd276909: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=40;
   mapp<=92;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=11795;
 end   
19'd276910: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=27;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=16592;
 end   
19'd276911: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=80;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=14976;
 end   
19'd276912: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=31;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=17374;
 end   
19'd276913: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=90;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=12872;
 end   
19'd276914: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=17;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd276915: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd277057: begin  
rid<=1;
end
19'd277058: begin  
end
19'd277059: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd277060: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd277061: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd277062: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd277063: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd277064: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd277065: begin  
rid<=0;
end
19'd277201: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=31;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=14574;
 end   
19'd277202: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=53;
   mapp<=26;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=16835;
 end   
19'd277203: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=71;
   mapp<=50;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=21216;
 end   
19'd277204: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=26;
   mapp<=77;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=14914;
 end   
19'd277205: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=91;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd277206: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=80;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd277207: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=20;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd277208: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=17;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd277209: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=53;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd277210: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=41;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd277211: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=74;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=34382;
 end   
19'd277212: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=22;
   mapp<=66;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=31177;
 end   
19'd277213: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=30;
   mapp<=47;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=37222;
 end   
19'd277214: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=39;
   mapp<=53;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=34684;
 end   
19'd277215: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=21;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd277216: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=68;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd277217: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=87;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd277218: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=7;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd277219: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=4;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd277220: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=95;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd277221: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd277363: begin  
rid<=1;
end
19'd277364: begin  
end
19'd277365: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd277366: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd277367: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd277368: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd277369: begin  
rid<=0;
end
19'd277501: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=21;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12050;
 end   
19'd277502: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=18;
   mapp<=37;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11732;
 end   
19'd277503: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=85;
   mapp<=48;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=14802;
 end   
19'd277504: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=37;
   mapp<=41;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=13634;
 end   
19'd277505: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=59;
   mapp<=81;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=15345;
 end   
19'd277506: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=61;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=13566;
 end   
19'd277507: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=66;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=14604;
 end   
19'd277508: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd277509: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd277510: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd277511: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd277512: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=96;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=24958;
 end   
19'd277513: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=30;
   mapp<=4;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=22401;
 end   
19'd277514: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=91;
   mapp<=2;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=28797;
 end   
19'd277515: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=98;
   mapp<=33;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=30137;
 end   
19'd277516: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=76;
   mapp<=45;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=34002;
 end   
19'd277517: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=37;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=34739;
 end   
19'd277518: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=67;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=41889;
 end   
19'd277519: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd277520: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd277521: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd277522: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd277523: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd277665: begin  
rid<=1;
end
19'd277666: begin  
end
19'd277667: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd277668: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd277669: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd277670: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd277671: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd277672: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd277673: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd277674: begin  
rid<=0;
end
19'd277801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=9;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9937;
 end   
19'd277802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=35;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=13585;
 end   
19'd277803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=26;
   mapp<=41;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9827;
 end   
19'd277804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=23;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd277805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=14;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd277806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=61;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd277807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=61;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd277808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=6;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd277809: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=20435;
 end   
19'd277810: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=92;
   mapp<=24;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=21770;
 end   
19'd277811: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=70;
   mapp<=55;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=14088;
 end   
19'd277812: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=94;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd277813: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=7;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd277814: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd277815: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=3;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd277816: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=76;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd277817: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd277959: begin  
rid<=1;
end
19'd277960: begin  
end
19'd277961: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd277962: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd277963: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd277964: begin  
rid<=0;
end
19'd278101: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=25;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8233;
 end   
19'd278102: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=89;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8523;
 end   
19'd278103: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=28;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7032;
 end   
19'd278104: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=69;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=9315;
 end   
19'd278105: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=59;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=7659;
 end   
19'd278106: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=46;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=9096;
 end   
19'd278107: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=79;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd278108: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=39;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=9595;
 end   
19'd278109: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=14;
   mapp<=36;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=11063;
 end   
19'd278110: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=62;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=10232;
 end   
19'd278111: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=51;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=11157;
 end   
19'd278112: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=20;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=11483;
 end   
19'd278113: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=94;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=11452;
 end   
19'd278114: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=8;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd278115: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd278257: begin  
rid<=1;
end
19'd278258: begin  
end
19'd278259: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd278260: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd278261: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd278262: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd278263: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd278264: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd278265: begin  
rid<=0;
end
19'd278401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=66;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4772;
 end   
19'd278402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=51;
   mapp<=28;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3012;
 end   
19'd278403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=88;
   mapp<=14;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9647;
 end   
19'd278404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=5;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7456;
 end   
19'd278405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=96;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=14867;
 end   
19'd278406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=25;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=13010;
 end   
19'd278407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=82;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=10219;
 end   
19'd278408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=81;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=8589;
 end   
19'd278409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=7;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=8862;
 end   
19'd278410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd278411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd278412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=74;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=14298;
 end   
19'd278413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=38;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=7744;
 end   
19'd278414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=40;
   mapp<=55;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=14157;
 end   
19'd278415: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=48;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=12408;
 end   
19'd278416: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=11;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=15801;
 end   
19'd278417: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=35;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=19040;
 end   
19'd278418: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=3;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=12601;
 end   
19'd278419: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=86;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=16553;
 end   
19'd278420: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=54;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=15298;
 end   
19'd278421: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd278422: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd278423: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd278565: begin  
rid<=1;
end
19'd278566: begin  
end
19'd278567: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd278568: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd278569: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd278570: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd278571: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd278572: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd278573: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd278574: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd278575: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd278576: begin  
rid<=0;
end
19'd278701: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=78;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=15615;
 end   
19'd278702: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=48;
   mapp<=37;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11786;
 end   
19'd278703: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=61;
   mapp<=83;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=14007;
 end   
19'd278704: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=44;
   mapp<=47;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=13214;
 end   
19'd278705: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=37;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=10472;
 end   
19'd278706: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=86;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=15462;
 end   
19'd278707: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=19;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=12561;
 end   
19'd278708: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=53;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd278709: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd278710: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=80;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd278711: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=4;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=24427;
 end   
19'd278712: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=30;
   mapp<=87;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=24510;
 end   
19'd278713: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=78;
   mapp<=69;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=25101;
 end   
19'd278714: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=52;
   mapp<=10;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=18321;
 end   
19'd278715: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=10;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=13250;
 end   
19'd278716: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=3;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=23131;
 end   
19'd278717: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=13;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=23914;
 end   
19'd278718: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=87;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd278719: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=31;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd278720: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=67;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd278721: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd278863: begin  
rid<=1;
end
19'd278864: begin  
end
19'd278865: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd278866: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd278867: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd278868: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd278869: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd278870: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd278871: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd278872: begin  
rid<=0;
end
19'd279001: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=2;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9685;
 end   
19'd279002: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=63;
   mapp<=16;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=20030;
 end   
19'd279003: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=13;
   mapp<=52;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=16122;
 end   
19'd279004: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=94;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd279005: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=56;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd279006: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=42;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd279007: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=85;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd279008: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=50;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd279009: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=93;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd279010: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=70;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=33670;
 end   
19'd279011: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=38;
   mapp<=73;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=41790;
 end   
19'd279012: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=81;
   mapp<=13;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=40024;
 end   
19'd279013: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=49;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd279014: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=99;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd279015: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=93;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd279016: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=95;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd279017: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=21;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd279018: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=92;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd279019: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd279161: begin  
rid<=1;
end
19'd279162: begin  
end
19'd279163: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd279164: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd279165: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd279166: begin  
rid<=0;
end
19'd279301: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=97;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7942;
 end   
19'd279302: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=48;
   mapp<=64;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9738;
 end   
19'd279303: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=54;
   mapp<=65;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11094;
 end   
19'd279304: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=4;
   mapp<=89;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=11096;
 end   
19'd279305: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=56;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd279306: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=76;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd279307: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=18;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd279308: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=84;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd279309: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=89;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=21103;
 end   
19'd279310: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=67;
   mapp<=98;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=19315;
 end   
19'd279311: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=21;
   mapp<=14;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=18997;
 end   
19'd279312: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=5;
   mapp<=48;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=18469;
 end   
19'd279313: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=6;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd279314: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=61;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd279315: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=66;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd279316: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=53;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd279317: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd279459: begin  
rid<=1;
end
19'd279460: begin  
end
19'd279461: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd279462: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd279463: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd279464: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd279465: begin  
rid<=0;
end
19'd279601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=17;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=19126;
 end   
19'd279602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=20;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=18575;
 end   
19'd279603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=1;
   mapp<=31;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=20058;
 end   
19'd279604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=39;
   mapp<=60;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=25593;
 end   
19'd279605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=57;
   mapp<=28;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=26631;
 end   
19'd279606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=90;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd279607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=74;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd279608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=50;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd279609: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=66;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd279610: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=95;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd279611: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=59;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd279612: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=40;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=37171;
 end   
19'd279613: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=39;
   mapp<=15;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=39464;
 end   
19'd279614: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=45;
   mapp<=94;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=43376;
 end   
19'd279615: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=72;
   mapp<=17;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=48827;
 end   
19'd279616: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=80;
   mapp<=26;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=51146;
 end   
19'd279617: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=38;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd279618: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=72;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd279619: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=50;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd279620: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=90;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd279621: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=67;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd279622: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=51;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd279623: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd279765: begin  
rid<=1;
end
19'd279766: begin  
end
19'd279767: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd279768: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd279769: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd279770: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd279771: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd279772: begin  
rid<=0;
end
19'd279901: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=77;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13375;
 end   
19'd279902: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=13;
   mapp<=8;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9126;
 end   
19'd279903: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=53;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd279904: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=51;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd279905: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=84;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd279906: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=68;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd279907: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=48;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17931;
 end   
19'd279908: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=88;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=14304;
 end   
19'd279909: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=95;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd279910: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=39;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd279911: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=15;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd279912: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=6;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd279913: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd280055: begin  
rid<=1;
end
19'd280056: begin  
end
19'd280057: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd280058: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd280059: begin  
rid<=0;
end
19'd280201: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=21;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11015;
 end   
19'd280202: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=47;
   mapp<=38;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12103;
 end   
19'd280203: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=58;
   mapp<=83;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=13482;
 end   
19'd280204: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=54;
   mapp<=55;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=15396;
 end   
19'd280205: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=40;
   mapp<=2;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=16301;
 end   
19'd280206: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=76;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd280207: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd280208: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd280209: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd280210: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=11;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=31071;
 end   
19'd280211: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=87;
   mapp<=98;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=35283;
 end   
19'd280212: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=88;
   mapp<=95;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=32903;
 end   
19'd280213: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=81;
   mapp<=11;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=26296;
 end   
19'd280214: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=38;
   mapp<=40;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=25573;
 end   
19'd280215: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=11;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd280216: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=42;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd280217: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=2;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd280218: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=39;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd280219: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd280361: begin  
rid<=1;
end
19'd280362: begin  
end
19'd280363: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd280364: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd280365: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd280366: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd280367: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd280368: begin  
rid<=0;
end
19'd280501: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=77;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11504;
 end   
19'd280502: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=32;
   mapp<=12;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9465;
 end   
19'd280503: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=47;
   mapp<=8;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8672;
 end   
19'd280504: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=8;
   mapp<=70;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=12543;
 end   
19'd280505: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=51;
   mapp<=94;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=15453;
 end   
19'd280506: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=83;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=11976;
 end   
19'd280507: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd280508: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd280509: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd280510: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd280511: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=72;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=27759;
 end   
19'd280512: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=28;
   mapp<=58;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=25897;
 end   
19'd280513: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=85;
   mapp<=68;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=24837;
 end   
19'd280514: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=61;
   mapp<=31;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=24196;
 end   
19'd280515: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=48;
   mapp<=73;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=27626;
 end   
19'd280516: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=68;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=23978;
 end   
19'd280517: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd280518: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd280519: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd280520: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd280521: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd280663: begin  
rid<=1;
end
19'd280664: begin  
end
19'd280665: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd280666: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd280667: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd280668: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd280669: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd280670: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd280671: begin  
rid<=0;
end
19'd280801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=26;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5789;
 end   
19'd280802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=53;
   mapp<=4;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11975;
 end   
19'd280803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=28;
   mapp<=7;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=13453;
 end   
19'd280804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=93;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd280805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=91;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd280806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd280807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd280808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=41;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=22179;
 end   
19'd280809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=63;
   mapp<=94;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=28627;
 end   
19'd280810: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=81;
   mapp<=92;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=24175;
 end   
19'd280811: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=13;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd280812: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=22;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd280813: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd280814: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd280815: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd280957: begin  
rid<=1;
end
19'd280958: begin  
end
19'd280959: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd280960: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd280961: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd280962: begin  
rid<=0;
end
19'd281101: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=36;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=25338;
 end   
19'd281102: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=10;
   mapp<=44;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=27091;
 end   
19'd281103: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=62;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd281104: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=91;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd281105: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=57;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd281106: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=55;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd281107: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=80;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd281108: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=59;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd281109: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=39;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd281110: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=26;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd281111: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=83;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=70685;
 end   
19'd281112: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=66;
   mapp<=90;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=67495;
 end   
19'd281113: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=44;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd281114: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=59;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd281115: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=93;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd281116: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=98;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd281117: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=25;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd281118: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=67;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd281119: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=65;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd281120: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=46;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd281121: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd281263: begin  
rid<=1;
end
19'd281264: begin  
end
19'd281265: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd281266: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd281267: begin  
rid<=0;
end
19'd281401: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=13;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6391;
 end   
19'd281402: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=7;
   mapp<=78;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2834;
 end   
19'd281403: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=76;
   mapp<=74;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5889;
 end   
19'd281404: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=17;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7608;
 end   
19'd281405: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=63;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4460;
 end   
19'd281406: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=91;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=8194;
 end   
19'd281407: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=39;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=5895;
 end   
19'd281408: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=88;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=2484;
 end   
19'd281409: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd281410: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd281411: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=4;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17989;
 end   
19'd281412: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=77;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=11368;
 end   
19'd281413: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=77;
   mapp<=57;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=14125;
 end   
19'd281414: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=49;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=16505;
 end   
19'd281415: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=55;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=10763;
 end   
19'd281416: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=58;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=10736;
 end   
19'd281417: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=21;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=11061;
 end   
19'd281418: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=9;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=13608;
 end   
19'd281419: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd281420: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd281421: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd281563: begin  
rid<=1;
end
19'd281564: begin  
end
19'd281565: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd281566: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd281567: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd281568: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd281569: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd281570: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd281571: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd281572: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd281573: begin  
rid<=0;
end
19'd281701: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=4;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=18438;
 end   
19'd281702: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=7;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd281703: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=29;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd281704: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=88;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd281705: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=78;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd281706: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=55;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd281707: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=69;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=37876;
 end   
19'd281708: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=73;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd281709: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=26;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd281710: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=89;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd281711: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=78;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd281712: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=6;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd281713: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd281855: begin  
rid<=1;
end
19'd281856: begin  
end
19'd281857: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd281858: begin  
rid<=0;
end
19'd282001: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=82;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=17935;
 end   
19'd282002: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=28;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd282003: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=68;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd282004: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd282005: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=80;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd282006: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=51;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd282007: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=18;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd282008: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=76;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd282009: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=53;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=27008;
 end   
19'd282010: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=39;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd282011: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=74;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd282012: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=6;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd282013: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=4;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd282014: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=28;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd282015: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=42;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd282016: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=83;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd282017: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd282159: begin  
rid<=1;
end
19'd282160: begin  
end
19'd282161: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd282162: begin  
rid<=0;
end
19'd282301: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=59;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1121;
 end   
19'd282302: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=63;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1207;
 end   
19'd282303: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=5;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=1321;
 end   
19'd282304: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=61;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=3647;
 end   
19'd282305: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd282447: begin  
rid<=1;
end
19'd282448: begin  
end
19'd282449: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd282450: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd282451: begin  
rid<=0;
end
19'd282601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=37;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1127;
 end   
19'd282602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=18;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1978;
 end   
19'd282603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=2;
   mapp<=2;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1650;
 end   
19'd282604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=78;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4316;
 end   
19'd282605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=76;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=3268;
 end   
19'd282606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd282607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd282608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=52;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=9900;
 end   
19'd282609: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=12;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=4636;
 end   
19'd282610: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=53;
   mapp<=89;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=8493;
 end   
19'd282611: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=30;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=11331;
 end   
19'd282612: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=35;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=10097;
 end   
19'd282613: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd282614: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd282615: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd282757: begin  
rid<=1;
end
19'd282758: begin  
end
19'd282759: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd282760: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd282761: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd282762: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd282763: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd282764: begin  
rid<=0;
end
19'd282901: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=13;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=19365;
 end   
19'd282902: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=81;
   mapp<=43;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=21821;
 end   
19'd282903: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=2;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd282904: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=54;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd282905: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=55;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd282906: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=58;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd282907: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=98;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd282908: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=76;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd282909: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=11;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd282910: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=42;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd282911: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=29;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=31417;
 end   
19'd282912: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=85;
   mapp<=28;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=36546;
 end   
19'd282913: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd282914: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=14;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd282915: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=14;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd282916: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=70;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd282917: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=25;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd282918: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=21;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd282919: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=6;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd282920: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=65;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd282921: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd283063: begin  
rid<=1;
end
19'd283064: begin  
end
19'd283065: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd283066: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd283067: begin  
rid<=0;
end
19'd283201: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=79;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5214;
 end   
19'd283202: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=25;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1985;
 end   
19'd283203: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=31;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2469;
 end   
19'd283204: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=39;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3111;
 end   
19'd283205: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=75;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5965;
 end   
19'd283206: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=55;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=4395;
 end   
19'd283207: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=32;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=2588;
 end   
19'd283208: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=89;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5392;
 end   
19'd283209: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=33;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=4922;
 end   
19'd283210: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=48;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=6741;
 end   
19'd283211: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=67;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=9074;
 end   
19'd283212: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=58;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=11127;
 end   
19'd283213: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=7;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=5018;
 end   
19'd283214: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=40;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=6148;
 end   
19'd283215: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd283357: begin  
rid<=1;
end
19'd283358: begin  
end
19'd283359: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd283360: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd283361: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd283362: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd283363: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd283364: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd283365: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd283366: begin  
rid<=0;
end
19'd283501: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=52;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=20454;
 end   
19'd283502: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=76;
   mapp<=47;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=18802;
 end   
19'd283503: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=95;
   mapp<=73;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=16979;
 end   
19'd283504: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=98;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd283505: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=87;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd283506: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=86;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd283507: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=68;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd283508: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=25;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd283509: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd283510: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=9;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd283511: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=68;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=41826;
 end   
19'd283512: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=78;
   mapp<=30;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=36155;
 end   
19'd283513: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=31;
   mapp<=75;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=30470;
 end   
19'd283514: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=61;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd283515: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=41;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd283516: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=15;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd283517: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=79;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd283518: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=39;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd283519: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=10;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd283520: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=92;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd283521: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd283663: begin  
rid<=1;
end
19'd283664: begin  
end
19'd283665: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd283666: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd283667: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd283668: begin  
rid<=0;
end
19'd283801: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=53;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4446;
 end   
19'd283802: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=52;
   mapp<=30;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6413;
 end   
19'd283803: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=67;
   mapp<=32;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6840;
 end   
19'd283804: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=47;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=8353;
 end   
19'd283805: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=40;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5608;
 end   
19'd283806: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=56;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=7655;
 end   
19'd283807: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=8;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=4028;
 end   
19'd283808: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=63;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=3818;
 end   
19'd283809: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=4;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=1989;
 end   
19'd283810: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd283811: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd283812: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=5;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=10431;
 end   
19'd283813: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=56;
   mapp<=99;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8859;
 end   
19'd283814: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=17;
   mapp<=23;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=9462;
 end   
19'd283815: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=39;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=10683;
 end   
19'd283816: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=19;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=10557;
 end   
19'd283817: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=63;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=13375;
 end   
19'd283818: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=78;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=8446;
 end   
19'd283819: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=61;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=7176;
 end   
19'd283820: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=36;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=6367;
 end   
19'd283821: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd283822: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd283823: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd283965: begin  
rid<=1;
end
19'd283966: begin  
end
19'd283967: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd283968: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd283969: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd283970: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd283971: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd283972: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd283973: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd283974: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd283975: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd283976: begin  
rid<=0;
end
19'd284101: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=33;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1815;
 end   
19'd284102: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=52;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2870;
 end   
19'd284103: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=24;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1340;
 end   
19'd284104: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=62;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3440;
 end   
19'd284105: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=39;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=2185;
 end   
19'd284106: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=18;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=2751;
 end   
19'd284107: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=12;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=3494;
 end   
19'd284108: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=25;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=2640;
 end   
19'd284109: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=56;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6352;
 end   
19'd284110: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=3;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=2341;
 end   
19'd284111: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd284253: begin  
rid<=1;
end
19'd284254: begin  
end
19'd284255: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd284256: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd284257: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd284258: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd284259: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd284260: begin  
rid<=0;
end
19'd284401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=64;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=20008;
 end   
19'd284402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=61;
   mapp<=31;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=18534;
 end   
19'd284403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=72;
   mapp<=73;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=15714;
 end   
19'd284404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=67;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd284405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=83;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd284406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=93;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd284407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=44;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd284408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=10;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd284409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=10;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd284410: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=30;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd284411: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=21;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=34340;
 end   
19'd284412: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=28;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=33332;
 end   
19'd284413: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=41;
   mapp<=9;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=32422;
 end   
19'd284414: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=92;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd284415: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=29;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd284416: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=93;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd284417: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=67;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd284418: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=25;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd284419: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=77;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd284420: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=48;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd284421: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd284563: begin  
rid<=1;
end
19'd284564: begin  
end
19'd284565: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd284566: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd284567: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd284568: begin  
rid<=0;
end
19'd284701: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=91;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16121;
 end   
19'd284702: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=25;
   mapp<=20;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=9825;
 end   
19'd284703: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=40;
   mapp<=17;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12694;
 end   
19'd284704: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=54;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd284705: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=5;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd284706: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=58;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd284707: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd284708: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd284709: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=83;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=43223;
 end   
19'd284710: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=99;
   mapp<=78;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=36225;
 end   
19'd284711: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=67;
   mapp<=94;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=37109;
 end   
19'd284712: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=39;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd284713: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=82;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd284714: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=94;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd284715: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd284716: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd284717: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd284859: begin  
rid<=1;
end
19'd284860: begin  
end
19'd284861: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd284862: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd284863: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd284864: begin  
rid<=0;
end
19'd285001: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=26;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=5550;
 end   
19'd285002: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=17;
   mapp<=63;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=3753;
 end   
19'd285003: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=9;
   mapp<=55;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3282;
 end   
19'd285004: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=45;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd285005: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd285006: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd285007: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=56;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=18113;
 end   
19'd285008: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=10;
   mapp<=57;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=17963;
 end   
19'd285009: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=95;
   mapp<=73;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=21071;
 end   
19'd285010: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=41;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd285011: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd285012: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd285013: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd285155: begin  
rid<=1;
end
19'd285156: begin  
end
19'd285157: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd285158: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd285159: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd285160: begin  
rid<=0;
end
19'd285301: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=5;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3480;
 end   
19'd285302: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=40;
   mapp<=82;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7924;
 end   
19'd285303: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=77;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8676;
 end   
19'd285304: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=68;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=9474;
 end   
19'd285305: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=82;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=10700;
 end   
19'd285306: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=90;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=4716;
 end   
19'd285307: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=13;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=7140;
 end   
19'd285308: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=80;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd285309: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=72;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5274;
 end   
19'd285310: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=17;
   mapp<=42;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=8305;
 end   
19'd285311: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=3;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=11199;
 end   
19'd285312: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=59;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=13257;
 end   
19'd285313: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=69;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=11987;
 end   
19'd285314: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=6;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=5352;
 end   
19'd285315: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=13;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=10569;
 end   
19'd285316: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=77;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd285317: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd285459: begin  
rid<=1;
end
19'd285460: begin  
end
19'd285461: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd285462: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd285463: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd285464: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd285465: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd285466: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd285467: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd285468: begin  
rid<=0;
end
19'd285601: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=54;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=18972;
 end   
19'd285602: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=78;
   mapp<=87;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=16486;
 end   
19'd285603: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=96;
   mapp<=87;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=13862;
 end   
19'd285604: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd285605: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd285606: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=86;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=25138;
 end   
19'd285607: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=25;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=29393;
 end   
19'd285608: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=59;
   mapp<=17;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=17519;
 end   
19'd285609: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd285610: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd285611: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd285753: begin  
rid<=1;
end
19'd285754: begin  
end
19'd285755: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd285756: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd285757: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd285758: begin  
rid<=0;
end
19'd285901: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=24;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12118;
 end   
19'd285902: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=29;
   mapp<=79;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10689;
 end   
19'd285903: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=57;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd285904: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=88;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd285905: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=50;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd285906: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd285907: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=55;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=22483;
 end   
19'd285908: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=26;
   mapp<=41;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=16182;
 end   
19'd285909: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=9;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd285910: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=79;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd285911: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=24;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd285912: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd285913: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd286055: begin  
rid<=1;
end
19'd286056: begin  
end
19'd286057: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd286058: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd286059: begin  
rid<=0;
end
19'd286201: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=37;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13889;
 end   
19'd286202: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=72;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd286203: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=50;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd286204: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=33;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd286205: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=38;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd286206: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=74;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd286207: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=36;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=26150;
 end   
19'd286208: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=14;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd286209: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=18;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd286210: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=40;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd286211: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=9;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd286212: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=86;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd286213: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd286355: begin  
rid<=1;
end
19'd286356: begin  
end
19'd286357: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd286358: begin  
rid<=0;
end
19'd286501: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=25;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=8129;
 end   
19'd286502: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=76;
   mapp<=60;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8712;
 end   
19'd286503: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=13;
   mapp<=28;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7191;
 end   
19'd286504: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=36;
   mapp<=55;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=8214;
 end   
19'd286505: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=58;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=6996;
 end   
19'd286506: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=50;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6438;
 end   
19'd286507: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=28;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=6541;
 end   
19'd286508: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=6;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd286509: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd286510: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=67;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd286511: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=56;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=16074;
 end   
19'd286512: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=66;
   mapp<=90;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=19458;
 end   
19'd286513: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=49;
   mapp<=21;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=12668;
 end   
19'd286514: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=2;
   mapp<=68;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=22287;
 end   
19'd286515: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=78;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=18210;
 end   
19'd286516: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=43;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=22626;
 end   
19'd286517: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=90;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=20415;
 end   
19'd286518: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=63;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd286519: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=90;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd286520: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=73;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd286521: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd286663: begin  
rid<=1;
end
19'd286664: begin  
end
19'd286665: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd286666: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd286667: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd286668: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd286669: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd286670: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd286671: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd286672: begin  
rid<=0;
end
19'd286801: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=84;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=20066;
 end   
19'd286802: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=69;
   mapp<=15;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15609;
 end   
19'd286803: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=63;
   mapp<=75;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=19327;
 end   
19'd286804: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=71;
   mapp<=19;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=16419;
 end   
19'd286805: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=54;
   mapp<=87;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=18924;
 end   
19'd286806: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=37;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd286807: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd286808: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd286809: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd286810: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd286811: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=2;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=40192;
 end   
19'd286812: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=45;
   mapp<=30;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=33200;
 end   
19'd286813: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=9;
   mapp<=20;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=38043;
 end   
19'd286814: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=84;
   mapp<=93;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=35095;
 end   
19'd286815: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=90;
   mapp<=91;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=35679;
 end   
19'd286816: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=40;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd286817: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd286818: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd286819: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd286820: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd286821: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd286963: begin  
rid<=1;
end
19'd286964: begin  
end
19'd286965: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd286966: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd286967: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd286968: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd286969: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd286970: begin  
rid<=0;
end
19'd287101: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=97;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=24654;
 end   
19'd287102: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=97;
   mapp<=85;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=22183;
 end   
19'd287103: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=86;
   mapp<=75;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=22814;
 end   
19'd287104: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=7;
   mapp<=63;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=22692;
 end   
19'd287105: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=1;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd287106: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=11;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd287107: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd287108: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd287109: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd287110: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=30;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=35317;
 end   
19'd287111: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=77;
   mapp<=21;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=33017;
 end   
19'd287112: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=55;
   mapp<=10;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=36282;
 end   
19'd287113: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=61;
   mapp<=46;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=37680;
 end   
19'd287114: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=34;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd287115: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=34;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd287116: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd287117: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd287118: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd287119: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd287261: begin  
rid<=1;
end
19'd287262: begin  
end
19'd287263: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd287264: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd287265: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd287266: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd287267: begin  
rid<=0;
end
19'd287401: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=36;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=15193;
 end   
19'd287402: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=75;
   mapp<=19;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=16163;
 end   
19'd287403: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=95;
   mapp<=9;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=21298;
 end   
19'd287404: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=74;
   mapp<=79;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=20231;
 end   
19'd287405: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=12;
   mapp<=58;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=17672;
 end   
19'd287406: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=75;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd287407: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=92;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd287408: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=73;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd287409: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=75;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd287410: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=81;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd287411: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=75;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd287412: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=31;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=29626;
 end   
19'd287413: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=1;
   mapp<=53;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=33456;
 end   
19'd287414: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=72;
   mapp<=42;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=38413;
 end   
19'd287415: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=67;
   mapp<=79;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=39550;
 end   
19'd287416: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=91;
   mapp<=5;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=33497;
 end   
19'd287417: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=10;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd287418: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=74;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd287419: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd287420: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=36;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd287421: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=32;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd287422: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=11;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd287423: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd287565: begin  
rid<=1;
end
19'd287566: begin  
end
19'd287567: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd287568: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd287569: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd287570: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd287571: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd287572: begin  
rid<=0;
end
19'd287701: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=34;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9190;
 end   
19'd287702: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=23;
   mapp<=64;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12349;
 end   
19'd287703: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=52;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd287704: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=77;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd287705: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=39;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd287706: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=34;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=19716;
 end   
19'd287707: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=69;
   mapp<=28;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=24782;
 end   
19'd287708: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=96;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd287709: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=87;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd287710: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd287711: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd287853: begin  
rid<=1;
end
19'd287854: begin  
end
19'd287855: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd287856: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd287857: begin  
rid<=0;
end
19'd288001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=84;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=4383;
 end   
19'd288002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=87;
   mapp<=33;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8176;
 end   
19'd288003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=62;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9665;
 end   
19'd288004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=51;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4836;
 end   
19'd288005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd288006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=7;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=11670;
 end   
19'd288007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=86;
   mapp<=84;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=14526;
 end   
19'd288008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=67;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=17702;
 end   
19'd288009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=88;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6570;
 end   
19'd288010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd288011: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd288153: begin  
rid<=1;
end
19'd288154: begin  
end
19'd288155: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd288156: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd288157: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd288158: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd288159: begin  
rid<=0;
end
19'd288301: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=38;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7092;
 end   
19'd288302: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=89;
   mapp<=12;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11378;
 end   
19'd288303: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=57;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd288304: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=46;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd288305: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=86;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd288306: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=87;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=22598;
 end   
19'd288307: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=11;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20132;
 end   
19'd288308: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=79;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd288309: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=3;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd288310: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd288311: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd288453: begin  
rid<=1;
end
19'd288454: begin  
end
19'd288455: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd288456: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd288457: begin  
rid<=0;
end
19'd288601: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=97;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11998;
 end   
19'd288602: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=39;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd288603: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=66;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd288604: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=94;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd288605: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=61;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=19617;
 end   
19'd288606: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=87;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd288607: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=55;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd288608: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=16;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd288609: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd288751: begin  
rid<=1;
end
19'd288752: begin  
end
19'd288753: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd288754: begin  
rid<=0;
end
19'd288901: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=58;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=23520;
 end   
19'd288902: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=93;
   mapp<=49;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=24283;
 end   
19'd288903: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=46;
   mapp<=75;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=25705;
 end   
19'd288904: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=18;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd288905: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=24;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd288906: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=46;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd288907: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=69;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd288908: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=68;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd288909: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=99;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd288910: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd288911: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd288912: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=78;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=40597;
 end   
19'd288913: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=65;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=44592;
 end   
19'd288914: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=20;
   mapp<=7;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=48062;
 end   
19'd288915: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=18;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd288916: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=61;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd288917: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=60;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd288918: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=47;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd288919: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=89;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd288920: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=93;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd288921: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd288922: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd288923: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd289065: begin  
rid<=1;
end
19'd289066: begin  
end
19'd289067: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd289068: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd289069: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd289070: begin  
rid<=0;
end
19'd289201: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=52;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=9505;
 end   
19'd289202: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=71;
   mapp<=1;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7607;
 end   
19'd289203: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=79;
   mapp<=74;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8613;
 end   
19'd289204: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=29;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=9561;
 end   
19'd289205: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=34;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=8745;
 end   
19'd289206: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=71;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=12398;
 end   
19'd289207: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd289208: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd289209: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=52;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=24569;
 end   
19'd289210: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=72;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=18463;
 end   
19'd289211: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=60;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=19513;
 end   
19'd289212: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=25;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=22273;
 end   
19'd289213: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=91;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=21469;
 end   
19'd289214: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=81;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=24122;
 end   
19'd289215: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd289216: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd289217: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd289359: begin  
rid<=1;
end
19'd289360: begin  
end
19'd289361: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd289362: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd289363: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd289364: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd289365: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd289366: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd289367: begin  
rid<=0;
end
19'd289501: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=78;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10883;
 end   
19'd289502: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=93;
   mapp<=70;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7053;
 end   
19'd289503: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=29;
   mapp<=19;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3767;
 end   
19'd289504: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=24;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=5258;
 end   
19'd289505: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=34;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=9500;
 end   
19'd289506: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=88;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=11750;
 end   
19'd289507: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=86;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=9599;
 end   
19'd289508: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=72;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=4857;
 end   
19'd289509: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=15;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd289510: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=11;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd289511: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=34;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=21592;
 end   
19'd289512: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=59;
   mapp<=76;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=16731;
 end   
19'd289513: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=81;
   mapp<=63;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=13443;
 end   
19'd289514: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=25;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=17531;
 end   
19'd289515: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=81;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=19124;
 end   
19'd289516: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=84;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=20624;
 end   
19'd289517: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=9;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=19330;
 end   
19'd289518: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=86;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=15538;
 end   
19'd289519: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=46;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd289520: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=69;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd289521: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd289663: begin  
rid<=1;
end
19'd289664: begin  
end
19'd289665: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd289666: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd289667: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd289668: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd289669: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd289670: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd289671: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd289672: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd289673: begin  
rid<=0;
end
19'd289801: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=96;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6528;
 end   
19'd289802: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=40;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2730;
 end   
19'd289803: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=20;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1380;
 end   
19'd289804: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=3;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=234;
 end   
19'd289805: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=19;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=1332;
 end   
19'd289806: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=5;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=390;
 end   
19'd289807: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=10;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=740;
 end   
19'd289808: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=88;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=6054;
 end   
19'd289809: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=67;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=4636;
 end   
19'd289810: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=42;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=2946;
 end   
19'd289811: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=45;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=8553;
 end   
19'd289812: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=46;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=4800;
 end   
19'd289813: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=60;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=4080;
 end   
19'd289814: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=48;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=2394;
 end   
19'd289815: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=76;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=4752;
 end   
19'd289816: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=14;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=1020;
 end   
19'd289817: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=80;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=4340;
 end   
19'd289818: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=54;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=8484;
 end   
19'd289819: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=93;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=8821;
 end   
19'd289820: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=51;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=5241;
 end   
19'd289821: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd289963: begin  
rid<=1;
end
19'd289964: begin  
end
19'd289965: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd289966: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd289967: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd289968: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd289969: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd289970: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd289971: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd289972: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd289973: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd289974: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd289975: begin  
rid<=0;
end
19'd290101: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=72;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=21273;
 end   
19'd290102: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=92;
   mapp<=79;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=16089;
 end   
19'd290103: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=8;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd290104: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=69;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd290105: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=5;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd290106: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=88;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd290107: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=44;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd290108: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd290109: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=11;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=38142;
 end   
19'd290110: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=70;
   mapp<=4;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=35906;
 end   
19'd290111: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=18;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd290112: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=50;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd290113: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=76;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd290114: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=69;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd290115: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=48;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd290116: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd290117: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd290259: begin  
rid<=1;
end
19'd290260: begin  
end
19'd290261: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd290262: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd290263: begin  
rid<=0;
end
19'd290401: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=15;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=20136;
 end   
19'd290402: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=70;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15546;
 end   
19'd290403: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=26;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd290404: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=9;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd290405: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=70;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd290406: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=78;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd290407: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=88;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd290408: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=23;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd290409: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd290410: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=3;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=39707;
 end   
19'd290411: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=38;
   mapp<=96;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=34483;
 end   
19'd290412: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=66;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd290413: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=36;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd290414: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=97;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd290415: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=81;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd290416: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=18;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd290417: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=40;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd290418: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd290419: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd290561: begin  
rid<=1;
end
19'd290562: begin  
end
19'd290563: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd290564: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd290565: begin  
rid<=0;
end
19'd290701: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=34;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=21256;
 end   
19'd290702: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=7;
   mapp<=26;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15335;
 end   
19'd290703: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=5;
   mapp<=85;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=19637;
 end   
19'd290704: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=62;
   mapp<=84;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=18807;
 end   
19'd290705: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=33;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd290706: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=34;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd290707: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=8;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd290708: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=91;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd290709: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=30;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd290710: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=81;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd290711: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=3;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd290712: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=78;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=51286;
 end   
19'd290713: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=1;
   mapp<=98;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=46620;
 end   
19'd290714: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=86;
   mapp<=72;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=53802;
 end   
19'd290715: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=19;
   mapp<=90;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=52005;
 end   
19'd290716: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=75;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd290717: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=67;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd290718: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=92;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd290719: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=51;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd290720: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=97;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd290721: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=15;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd290722: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=57;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd290723: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd290865: begin  
rid<=1;
end
19'd290866: begin  
end
19'd290867: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd290868: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd290869: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd290870: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd290871: begin  
rid<=0;
end
19'd291001: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=7;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1216;
 end   
19'd291002: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=24;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd291003: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=25;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=4116;
 end   
19'd291004: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=80;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd291005: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd291147: begin  
rid<=1;
end
19'd291148: begin  
end
19'd291149: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd291150: begin  
rid<=0;
end
19'd291301: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=71;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1846;
 end   
19'd291302: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=23;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1643;
 end   
19'd291303: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=4;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=304;
 end   
19'd291304: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=57;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4077;
 end   
19'd291305: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=5;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=395;
 end   
19'd291306: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=96;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6866;
 end   
19'd291307: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=5;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=415;
 end   
19'd291308: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=33;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=2413;
 end   
19'd291309: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=36;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=2818;
 end   
19'd291310: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=27;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=2615;
 end   
19'd291311: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=2824;
 end   
19'd291312: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=8;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=4365;
 end   
19'd291313: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=82;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=3347;
 end   
19'd291314: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=17;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=7478;
 end   
19'd291315: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=64;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=2719;
 end   
19'd291316: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=10;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=2773;
 end   
19'd291317: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd291459: begin  
rid<=1;
end
19'd291460: begin  
end
19'd291461: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd291462: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd291463: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd291464: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd291465: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd291466: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd291467: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd291468: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd291469: begin  
rid<=0;
end
19'd291601: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=89;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13612;
 end   
19'd291602: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=55;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd291603: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=74;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd291604: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=46;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd291605: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=27;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=23906;
 end   
19'd291606: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=88;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd291607: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=15;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd291608: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=70;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd291609: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd291751: begin  
rid<=1;
end
19'd291752: begin  
end
19'd291753: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd291754: begin  
rid<=0;
end
19'd291901: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=93;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=18359;
 end   
19'd291902: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=11;
   mapp<=58;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12950;
 end   
19'd291903: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=17;
   mapp<=52;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=14536;
 end   
19'd291904: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=39;
   mapp<=97;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=20729;
 end   
19'd291905: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=92;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd291906: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=12;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd291907: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd291908: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd291909: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd291910: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=77;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=29231;
 end   
19'd291911: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=74;
   mapp<=41;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=21125;
 end   
19'd291912: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=30;
   mapp<=12;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=22092;
 end   
19'd291913: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=12;
   mapp<=6;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=28049;
 end   
19'd291914: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=62;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd291915: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=41;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd291916: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd291917: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd291918: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd291919: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd292061: begin  
rid<=1;
end
19'd292062: begin  
end
19'd292063: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd292064: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd292065: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd292066: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd292067: begin  
rid<=0;
end
19'd292201: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=7243;
 end   
19'd292202: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=31;
   mapp<=34;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10201;
 end   
19'd292203: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=60;
   mapp<=53;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=9842;
 end   
19'd292204: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=78;
   mapp<=32;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=7429;
 end   
19'd292205: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=9;
   mapp<=57;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=7964;
 end   
19'd292206: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=54;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=6284;
 end   
19'd292207: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=65;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd292208: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=9;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd292209: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd292210: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=21;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd292211: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=9;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=13879;
 end   
19'd292212: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=31;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=16089;
 end   
19'd292213: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=37;
   mapp<=77;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=19620;
 end   
19'd292214: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=9;
   mapp<=36;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=18777;
 end   
19'd292215: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=38;
   mapp<=55;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=24234;
 end   
19'd292216: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=28;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=19936;
 end   
19'd292217: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=79;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd292218: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=86;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd292219: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd292220: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=3;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd292221: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd292363: begin  
rid<=1;
end
19'd292364: begin  
end
19'd292365: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd292366: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd292367: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd292368: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd292369: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd292370: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd292371: begin  
rid<=0;
end
19'd292501: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=34;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6686;
 end   
19'd292502: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=82;
   mapp<=27;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8753;
 end   
19'd292503: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=38;
   mapp<=45;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8168;
 end   
19'd292504: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=32;
   mapp<=47;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6954;
 end   
19'd292505: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=69;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=5920;
 end   
19'd292506: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=59;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd292507: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=26;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd292508: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd292509: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=19;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=18065;
 end   
19'd292510: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=11;
   mapp<=43;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=23271;
 end   
19'd292511: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=73;
   mapp<=80;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=26923;
 end   
19'd292512: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=91;
   mapp<=35;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=23511;
 end   
19'd292513: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=86;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=23272;
 end   
19'd292514: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=21;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd292515: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd292516: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=85;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd292517: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd292659: begin  
rid<=1;
end
19'd292660: begin  
end
19'd292661: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd292662: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd292663: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd292664: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd292665: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd292666: begin  
rid<=0;
end
19'd292801: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=67;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11376;
 end   
19'd292802: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=29;
   mapp<=15;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=7498;
 end   
19'd292803: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=78;
   mapp<=81;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11586;
 end   
19'd292804: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=53;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=8646;
 end   
19'd292805: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=59;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=11324;
 end   
19'd292806: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=43;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=8937;
 end   
19'd292807: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=78;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=10500;
 end   
19'd292808: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd292809: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd292810: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=1;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=11613;
 end   
19'd292811: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=11;
   mapp<=21;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=10494;
 end   
19'd292812: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=85;
   mapp<=0;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=14776;
 end   
19'd292813: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=35;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=16949;
 end   
19'd292814: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=33;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=16970;
 end   
19'd292815: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=93;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=15659;
 end   
19'd292816: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=54;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=13970;
 end   
19'd292817: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd292818: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd292819: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd292961: begin  
rid<=1;
end
19'd292962: begin  
end
19'd292963: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd292964: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd292965: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd292966: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd292967: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd292968: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd292969: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd292970: begin  
rid<=0;
end
19'd293101: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=41;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=3593;
 end   
19'd293102: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=70;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6012;
 end   
19'd293103: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=67;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=3467;
 end   
19'd293104: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd293105: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=92;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=5192;
 end   
19'd293106: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=5;
   mapp<=7;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=7021;
 end   
19'd293107: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=73;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=10273;
 end   
19'd293108: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd293109: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd293251: begin  
rid<=1;
end
19'd293252: begin  
end
19'd293253: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd293254: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd293255: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd293256: begin  
rid<=0;
end
19'd293401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=14;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11675;
 end   
19'd293402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=44;
   mapp<=92;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11201;
 end   
19'd293403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=2;
   mapp<=38;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=11606;
 end   
19'd293404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=58;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd293405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=51;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd293406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=19;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd293407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=26;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd293408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=18;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd293409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=13;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd293410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd293411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd293412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=97;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=26754;
 end   
19'd293413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=21;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=34047;
 end   
19'd293414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=57;
   mapp<=40;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=36902;
 end   
19'd293415: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=6;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd293416: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=4;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd293417: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=72;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd293418: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=88;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd293419: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=20;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd293420: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=66;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd293421: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd293422: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd293423: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd293565: begin  
rid<=1;
end
19'd293566: begin  
end
19'd293567: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd293568: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd293569: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd293570: begin  
rid<=0;
end
19'd293701: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=11627;
 end   
19'd293702: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=26;
   mapp<=36;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15137;
 end   
19'd293703: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=78;
   mapp<=64;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=13880;
 end   
19'd293704: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=12;
   mapp<=99;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=14076;
 end   
19'd293705: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=89;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd293706: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=6;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd293707: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=76;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd293708: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=24;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd293709: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=14;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd293710: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=69;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd293711: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=52;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=38449;
 end   
19'd293712: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=95;
   mapp<=62;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=41955;
 end   
19'd293713: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=66;
   mapp<=73;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=39455;
 end   
19'd293714: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=90;
   mapp<=81;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=39409;
 end   
19'd293715: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=81;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd293716: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=20;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd293717: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=63;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd293718: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=84;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd293719: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=72;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd293720: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd293721: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd293863: begin  
rid<=1;
end
19'd293864: begin  
end
19'd293865: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd293866: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd293867: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd293868: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd293869: begin  
rid<=0;
end
19'd294001: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=24;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16246;
 end   
19'd294002: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=13;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd294003: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=45;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd294004: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=17;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd294005: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=62;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd294006: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=42;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd294007: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=59;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd294008: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=83;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd294009: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=25;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=48628;
 end   
19'd294010: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=4;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd294011: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=40;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd294012: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=76;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd294013: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=44;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd294014: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=82;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd294015: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=80;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd294016: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=80;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd294017: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd294159: begin  
rid<=1;
end
19'd294160: begin  
end
19'd294161: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd294162: begin  
rid<=0;
end
19'd294301: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=32;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=12518;
 end   
19'd294302: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=51;
   mapp<=98;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11949;
 end   
19'd294303: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=57;
   mapp<=16;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=16612;
 end   
19'd294304: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=91;
   mapp<=11;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=14219;
 end   
19'd294305: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=64;
   mapp<=72;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=9706;
 end   
19'd294306: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=35;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd294307: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd294308: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=64;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd294309: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=40;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd294310: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=44;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd294311: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=92;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=17744;
 end   
19'd294312: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=26;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=17430;
 end   
19'd294313: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=16;
   mapp<=50;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=21857;
 end   
19'd294314: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=70;
   mapp<=20;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=20743;
 end   
19'd294315: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=1;
   mapp<=25;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=17534;
 end   
19'd294316: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=21;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd294317: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd294318: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=39;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd294319: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=72;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd294320: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=83;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd294321: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd294463: begin  
rid<=1;
end
19'd294464: begin  
end
19'd294465: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd294466: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd294467: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd294468: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd294469: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd294470: begin  
rid<=0;
end
19'd294601: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=29;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6160;
 end   
19'd294602: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=71;
   mapp<=4;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=5475;
 end   
19'd294603: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=97;
   mapp<=33;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=7672;
 end   
19'd294604: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=76;
   mapp<=2;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6954;
 end   
19'd294605: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=37;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=8036;
 end   
19'd294606: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd294607: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd294608: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd294609: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=83;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=19275;
 end   
19'd294610: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=75;
   mapp<=89;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=17938;
 end   
19'd294611: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=17;
   mapp<=43;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=16336;
 end   
19'd294612: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=19;
   mapp<=34;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=16154;
 end   
19'd294613: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=67;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=20543;
 end   
19'd294614: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd294615: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd294616: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd294617: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd294759: begin  
rid<=1;
end
19'd294760: begin  
end
19'd294761: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd294762: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd294763: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd294764: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd294765: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd294766: begin  
rid<=0;
end
19'd294901: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=61;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10900;
 end   
19'd294902: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=95;
   mapp<=79;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8630;
 end   
19'd294903: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=1;
   mapp<=40;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=2620;
 end   
19'd294904: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=1;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=6309;
 end   
19'd294905: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd294906: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd294907: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd294908: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=91;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=22018;
 end   
19'd294909: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=19;
   mapp<=30;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=20244;
 end   
19'd294910: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=66;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=18365;
 end   
19'd294911: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=78;
   mapp<=27;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=16658;
 end   
19'd294912: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd294913: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd294914: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd294915: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd295057: begin  
rid<=1;
end
19'd295058: begin  
end
19'd295059: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd295060: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd295061: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd295062: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd295063: begin  
rid<=0;
end
19'd295201: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=53;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1855;
 end   
19'd295202: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=29;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=1025;
 end   
19'd295203: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=53;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=1875;
 end   
19'd295204: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=52;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=1850;
 end   
19'd295205: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=10;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=390;
 end   
19'd295206: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=58;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=2080;
 end   
19'd295207: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=37;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=2484;
 end   
19'd295208: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=13;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=1246;
 end   
19'd295209: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=34;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=2453;
 end   
19'd295210: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=51;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=2717;
 end   
19'd295211: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=93;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=1971;
 end   
19'd295212: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=28;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=2556;
 end   
19'd295213: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd295355: begin  
rid<=1;
end
19'd295356: begin  
end
19'd295357: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd295358: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd295359: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd295360: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd295361: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd295362: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd295363: begin  
rid<=0;
end
19'd295501: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=32;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=16934;
 end   
19'd295502: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=27;
   mapp<=9;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=14916;
 end   
19'd295503: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=32;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd295504: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=28;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd295505: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=82;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd295506: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=68;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd295507: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=65;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd295508: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=97;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd295509: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd295510: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=62;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=41747;
 end   
19'd295511: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=94;
   mapp<=18;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=38987;
 end   
19'd295512: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=17;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd295513: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=34;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd295514: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=29;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd295515: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=40;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd295516: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=86;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd295517: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=82;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd295518: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd295519: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd295661: begin  
rid<=1;
end
19'd295662: begin  
end
19'd295663: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd295664: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd295665: begin  
rid<=0;
end
19'd295801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=17;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=22722;
 end   
19'd295802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=63;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=20454;
 end   
19'd295803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=3;
   mapp<=76;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=25712;
 end   
19'd295804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=52;
   mapp<=61;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=28444;
 end   
19'd295805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=86;
   mapp<=66;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=27033;
 end   
19'd295806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=76;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd295807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=74;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd295808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=3;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd295809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=64;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd295810: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=80;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd295811: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=48;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd295812: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=72;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=43367;
 end   
19'd295813: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=53;
   mapp<=86;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=40553;
 end   
19'd295814: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=8;
   mapp<=65;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=47164;
 end   
19'd295815: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=82;
   mapp<=46;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=52538;
 end   
19'd295816: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=37;
   mapp<=63;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=52865;
 end   
19'd295817: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=94;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd295818: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=33;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd295819: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=22;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd295820: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=50;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd295821: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=54;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd295822: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=85;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd295823: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd295965: begin  
rid<=1;
end
19'd295966: begin  
end
19'd295967: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd295968: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd295969: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd295970: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd295971: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd295972: begin  
rid<=0;
end
19'd296101: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=39;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6695;
 end   
19'd296102: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=31;
   mapp<=43;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=12629;
 end   
19'd296103: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=17;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd296104: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=61;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd296105: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=11;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd296106: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=95;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd296107: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd296108: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=27;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=13744;
 end   
19'd296109: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=6;
   mapp<=79;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=23293;
 end   
19'd296110: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=55;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd296111: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=10;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd296112: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=78;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd296113: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=36;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd296114: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd296115: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd296257: begin  
rid<=1;
end
19'd296258: begin  
end
19'd296259: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd296260: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd296261: begin  
rid<=0;
end
19'd296401: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=59;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=28443;
 end   
19'd296402: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=45;
   mapp<=88;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=24389;
 end   
19'd296403: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=22;
   mapp<=97;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=20627;
 end   
19'd296404: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=10;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd296405: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=8;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd296406: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=55;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd296407: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=80;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd296408: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=74;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd296409: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=82;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd296410: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=33;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[9]<=0;
 end   
19'd296411: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=28;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[10]<=0;
 end   
19'd296412: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=37;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=46402;
 end   
19'd296413: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=33;
   mapp<=65;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=44127;
 end   
19'd296414: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=55;
   mapp<=62;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=43237;
 end   
19'd296415: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=17;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd296416: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=55;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd296417: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=92;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd296418: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=10;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd296419: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=27;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd296420: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=30;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd296421: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=77;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[9]<=0;
 end   
19'd296422: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=41;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[10]<=0;
 end   
19'd296423: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd296565: begin  
rid<=1;
end
19'd296566: begin  
end
19'd296567: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd296568: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd296569: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd296570: begin  
rid<=0;
end
19'd296701: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=48;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13068;
 end   
19'd296702: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=60;
   mapp<=62;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=10340;
 end   
19'd296703: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=43;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd296704: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=65;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd296705: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=0;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd296706: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=75;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=26380;
 end   
19'd296707: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=73;
   mapp<=73;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=22762;
 end   
19'd296708: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=8;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd296709: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=84;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd296710: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=0;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd296711: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd296853: begin  
rid<=1;
end
19'd296854: begin  
end
19'd296855: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd296856: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd296857: begin  
rid<=0;
end
19'd297001: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=28;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=2212;
 end   
19'd297002: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=0;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=4957;
 end   
19'd297003: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=51;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=6280;
 end   
19'd297004: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=23;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=3108;
 end   
19'd297005: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=13;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=4850;
 end   
19'd297006: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=39;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=3810;
 end   
19'd297007: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=7;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=7597;
 end   
19'd297008: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=72;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=7116;
 end   
19'd297009: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=14;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd297010: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=91;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=10925;
 end   
19'd297011: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=94;
   mapp<=53;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=11302;
 end   
19'd297012: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=47;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=9108;
 end   
19'd297013: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=17;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=6508;
 end   
19'd297014: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=51;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=11128;
 end   
19'd297015: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=79;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=11236;
 end   
19'd297016: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=79;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=13751;
 end   
19'd297017: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=55;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=9636;
 end   
19'd297018: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=5;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd297019: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd297161: begin  
rid<=1;
end
19'd297162: begin  
end
19'd297163: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd297164: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd297165: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd297166: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd297167: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd297168: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd297169: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd297170: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd297171: begin  
rid<=0;
end
19'd297301: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=81;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10146;
 end   
19'd297302: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=8;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[1]<=0;
 end   
19'd297303: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=9;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd297304: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=99;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd297305: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=46;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd297306: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=85;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=29845;
 end   
19'd297307: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=77;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[1]<=0;
 end   
19'd297308: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=80;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd297309: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=73;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd297310: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=67;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd297311: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd297453: begin  
rid<=1;
end
19'd297454: begin  
end
19'd297455: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd297456: begin  
rid<=0;
end
19'd297601: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=85;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=28464;
 end   
19'd297602: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=85;
   mapp<=76;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=19375;
 end   
19'd297603: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=30;
   mapp<=33;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=16372;
 end   
19'd297604: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=89;
   mapp<=92;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=20875;
 end   
19'd297605: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=34;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd297606: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=55;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd297607: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=19;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd297608: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd297609: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=93;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd297610: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=88;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=45993;
 end   
19'd297611: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=84;
   mapp<=38;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=34091;
 end   
19'd297612: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=97;
   mapp<=8;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=35531;
 end   
19'd297613: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=94;
   mapp<=20;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=40847;
 end   
19'd297614: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=47;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd297615: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=6;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd297616: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=28;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd297617: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=83;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd297618: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=55;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd297619: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd297761: begin  
rid<=1;
end
19'd297762: begin  
end
19'd297763: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd297764: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd297765: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd297766: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd297767: begin  
rid<=0;
end
19'd297901: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=96;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=13571;
 end   
19'd297902: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=37;
   mapp<=31;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=15181;
 end   
19'd297903: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=4;
   mapp<=58;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=15369;
 end   
19'd297904: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=78;
   mapp<=87;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=16422;
 end   
19'd297905: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=83;
   mapp<=42;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=17702;
 end   
19'd297906: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=61;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd297907: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=65;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd297908: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=73;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd297909: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=95;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[8]<=0;
 end   
19'd297910: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=11;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=28489;
 end   
19'd297911: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=29;
   mapp<=28;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=28005;
 end   
19'd297912: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=91;
   mapp<=79;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=30270;
 end   
19'd297913: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=59;
   mapp<=93;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=33032;
 end   
19'd297914: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=33;
   mapp<=24;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=35723;
 end   
19'd297915: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=36;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd297916: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=84;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd297917: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=67;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd297918: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=93;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[8]<=0;
 end   
19'd297919: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd298061: begin  
rid<=1;
end
19'd298062: begin  
end
19'd298063: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd298064: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd298065: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd298066: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd298067: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd298068: begin  
rid<=0;
end
19'd298201: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=21;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1764;
 end   
19'd298202: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=96;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=8074;
 end   
19'd298203: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=60;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=5060;
 end   
19'd298204: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=50;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=4230;
 end   
19'd298205: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=94;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=7936;
 end   
19'd298206: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=25;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=2150;
 end   
19'd298207: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=5;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=480;
 end   
19'd298208: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=1;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[7]<=154;
 end   
19'd298209: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=59;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[8]<=5036;
 end   
19'd298210: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=20;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[9]<=1770;
 end   
19'd298211: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=94;
   mapp<=0;
   pp<=100;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[10]<=7996;
 end   
19'd298212: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=15;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=2109;
 end   
19'd298213: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=89;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=10121;
 end   
19'd298214: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=67;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=6601;
 end   
19'd298215: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=40;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=5150;
 end   
19'd298216: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=86;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=9914;
 end   
19'd298217: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=12;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=2426;
 end   
19'd298218: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=16;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=848;
 end   
19'd298219: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=9;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[7]<=361;
 end   
19'd298220: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=40;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[8]<=5956;
 end   
19'd298221: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=42;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[9]<=2736;
 end   
19'd298222: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=60;
   mapp<=0;
   pp<=100;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[10]<=9376;
 end   
19'd298223: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd298365: begin  
rid<=1;
end
19'd298366: begin  
end
19'd298367: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd298368: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd298369: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd298370: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd298371: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd298372: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd298373: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd298374: begin  
check0<=expctdoutput[7]-outcheck0;
end
19'd298375: begin  
check0<=expctdoutput[8]-outcheck0;
end
19'd298376: begin  
check0<=expctdoutput[9]-outcheck0;
end
19'd298377: begin  
check0<=expctdoutput[10]-outcheck0;
end
19'd298378: begin  
rid<=0;
end
19'd298501: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=55;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=6742;
 end   
19'd298502: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=5;
   mapp<=42;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=6604;
 end   
19'd298503: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=41;
   mapp<=52;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=8628;
 end   
19'd298504: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=86;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=11572;
 end   
19'd298505: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=33;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd298506: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=63;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd298507: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=26;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=10897;
 end   
19'd298508: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=73;
   mapp<=19;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=13702;
 end   
19'd298509: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=31;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=16812;
 end   
19'd298510: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=69;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=18541;
 end   
19'd298511: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd298512: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=53;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd298513: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd298655: begin  
rid<=1;
end
19'd298656: begin  
end
19'd298657: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd298658: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd298659: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd298660: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd298661: begin  
rid<=0;
end
19'd298801: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=52;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=23272;
 end   
19'd298802: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=41;
   mapp<=80;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=27260;
 end   
19'd298803: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=69;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd298804: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=67;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd298805: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=69;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd298806: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=16;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[5]<=0;
 end   
19'd298807: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=73;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[6]<=0;
 end   
19'd298808: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[7]<=0;
 end   
19'd298809: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=90;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=42912;
 end   
19'd298810: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=90;
   mapp<=26;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=43268;
 end   
19'd298811: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=12;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd298812: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=55;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd298813: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=47;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd298814: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=36;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[5]<=0;
 end   
19'd298815: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=12;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[6]<=0;
 end   
19'd298816: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[7]<=0;
 end   
19'd298817: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd298959: begin  
rid<=1;
end
19'd298960: begin  
end
19'd298961: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd298962: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd298963: begin  
rid<=0;
end
19'd299101: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=36;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=10434;
 end   
19'd299102: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=89;
   mapp<=66;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=11921;
 end   
19'd299103: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=48;
   mapp<=71;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=12139;
 end   
19'd299104: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd299105: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=0;
 expctdoutput[4]<=0;
 end   
19'd299106: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=46;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=28778;
 end   
19'd299107: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=62;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=26513;
 end   
19'd299108: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=99;
   mapp<=92;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=23976;
 end   
19'd299109: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd299110: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
   idp<=1;
 expctdoutput[4]<=0;
 end   
19'd299111: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd299253: begin  
rid<=1;
end
19'd299254: begin  
end
19'd299255: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd299256: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd299257: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd299258: begin  
rid<=0;
end
19'd299401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=4;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1935;
 end   
19'd299402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=55;
   mapp<=13;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=2783;
 end   
19'd299403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=60;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[2]<=0;
 end   
19'd299404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=47;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=0;
 expctdoutput[3]<=0;
 end   
19'd299405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=54;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=15106;
 end   
19'd299406: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=71;
   mapp<=71;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=17121;
 end   
19'd299407: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=96;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[2]<=0;
 end   
19'd299408: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=17;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
   idp<=1;
 expctdoutput[3]<=0;
 end   
19'd299409: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd299551: begin  
rid<=1;
end
19'd299552: begin  
end
19'd299553: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd299554: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd299555: begin  
rid<=0;
end
19'd299701: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=38;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[0]<=1938;
 end   
19'd299702: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=5;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[1]<=265;
 end   
19'd299703: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=17;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[2]<=887;
 end   
19'd299704: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=48;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[3]<=2478;
 end   
19'd299705: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=17;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[4]<=907;
 end   
19'd299706: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=27;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[5]<=1427;
 end   
19'd299707: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=75;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=0;
 expctdoutput[6]<=3885;
 end   
19'd299708: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=21;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[0]<=2652;
 end   
19'd299709: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=34;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[1]<=1421;
 end   
19'd299710: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=24;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[2]<=1703;
 end   
19'd299711: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=70;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[3]<=4858;
 end   
19'd299712: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=14;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[4]<=1383;
 end   
19'd299713: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=2;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[5]<=1495;
 end   
19'd299714: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=8;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
   idp<=1;
 expctdoutput[6]<=4157;
 end   
19'd299715: begin  
   gm<=0;
   gf<=0;
   gp<=0;
end
19'd299857: begin  
rid<=1;
end
19'd299858: begin  
end
19'd299859: begin  
check0<=expctdoutput[0]-outcheck0;
end
19'd299860: begin  
check0<=expctdoutput[1]-outcheck0;
end
19'd299861: begin  
check0<=expctdoutput[2]-outcheck0;
end
19'd299862: begin  
check0<=expctdoutput[3]-outcheck0;
end
19'd299863: begin  
check0<=expctdoutput[4]-outcheck0;
end
19'd299864: begin  
check0<=expctdoutput[5]-outcheck0;
end
19'd299865: begin  
check0<=expctdoutput[6]-outcheck0;
end
19'd299866: begin  
rid<=0;
end


//XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXx



 endcase

end


endmodule

