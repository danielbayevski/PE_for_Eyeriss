`include "Eyeriss_PE.v"
`include "clock.sv"
`include "FIFObuffer16b_16b.v"
module Eyeriss_PE_tb();

reg [17:0] dismod;
reg clrr;
reg [15:0] filterp,mapp,pp;
reg gm, gf, gp;
wire [15:0] filter,map,p;
clock clk(.CLK(CLK));
wire [31:0] out, done;
reg [3:0]maplen;
reg [7:0] fillen;
reg [31:0] expctdoutput [11:0];
wire [15:0] psum_out;
wire clrrr;
assign clrrr=!clrr;
wire pnm;


Eyeriss_PE pe(.map(map), .filter(filter),.Psum_from_GLB(p),.Psum_from_PE(16'b0),.getdata_fil(gf),.getdata_map(gm),.getdata_psum(gp),
.id_in(8'b1),.stall(1'b0),.psum_i_empty(1'b0),.psum_i_full(1'b0),
 
.CLK(CLK),
.clr(~clr),
.conf_i({6'b110000,maplen,fillen,8'b00000001}),
							// enable, GLB input, 0 mult bit, 4 map len,7 fitler len, id =1; 
							//	1bit	1bit 	   4bit			4bit		8bit		8bit 
.ready(),.psum_out(psum_out),.psum_o_empty(pnm),.psum_o_full()
);
/*        conf_i = 
  wire conf_enable;                                               1
	wire conf_psum_input;  //0- psum from PE, 1-psum from GLB     1
    wire [3:0]mult_bit_select;                                    0000
	wire [3:0] conf_maplen;                                       0010
    wire [7:0] conf_filterlen;                                    00000011
	wire [7:0] conf_id;                                           00000001
	=> 11000000100000001100000001
*/                 
reg rid;
reg[15:0]check;
wire [15:0] outcheck;
assign clr=clrr;
assign filter=filterp;
assign map=mapp;
assign p=pp;
initial rid=0;
initial check=0;

FIFObuffer16b_16b Fifo_outside(
.Clk(CLK),
.dataIn(psum_out),
.RD(rid),
.WR(!pnm),
.EN(1'b1),
.dataOut(outcheck),
.Rst(clr),.EMPTY(), 
.FULL()
);

wire [15:0]testwire;
wire eme,emr,fle,flr;
reg wr;

/*
FIFObuffer16b_16b test_e(
.Clk(CLK),
.dataIn(dismod),
.RD(!flr),
.WR(wr),
.EN(1'b1),
.dataOut(testwire),
.Rst(clrr),.EMPTY(eme), 
.FULL(fle)
);

FIFObuffer16b_16b test_r(
.Clk(CLK),
.dataIn(testwire),
.RD(1'b0),
.WR(!eme),
.EN(1'b1),
.dataOut(),
.Rst(clrr),.EMPTY(emr), 
.FULL(flr)
);
*/

 

//TODO: more tests,how about a test every 1000 CLKS 
	
 initial dismod=0;
always@(posedge CLK) begin
 dismod<=dismod+1;
 
 case(dismod)
/* 
 default: 
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
   clrr<=0;
   filterp<=0;
   mapp<=0;
   
   end 
 */
//XXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXXX

18'd0: begin
clrr<=1;  
 end   
18'd1: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=45;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=21977;
 end   
18'd2: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=81;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=23436;
 end   
18'd3: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=27;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd4: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=61;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd5: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=91;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd6: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=95;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd7: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=42;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd8: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=27;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd9: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=36;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd10: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=91;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd11: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd12: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd13: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21977;
 end   
18'd14: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21977;
 end   
18'd15: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21977;
 end   
18'd16: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21977;
 end   
18'd17: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21977;
 end   
18'd18: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21977;
 end   
18'd19: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21977;
 end   
18'd142: begin  
rid<=1;
end
18'd143: begin  
end
18'd144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd146: begin  
rid<=0;
end
18'd201: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=26;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=24923;
 end   
18'd202: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=71;
   mapp<=92;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=23776;
 end   
18'd203: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=38;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd204: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=69;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd205: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=12;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd206: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=67;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd207: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=99;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd208: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=35;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd209: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=94;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd210: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd211: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd212: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd213: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24923;
 end   
18'd214: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24923;
 end   
18'd215: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24923;
 end   
18'd216: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24923;
 end   
18'd217: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24923;
 end   
18'd342: begin  
rid<=1;
end
18'd343: begin  
end
18'd344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd346: begin  
rid<=0;
end
18'd401: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=11;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11767;
 end   
18'd402: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=53;
   mapp<=33;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=12209;
 end   
18'd403: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=68;
   mapp<=73;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12584;
 end   
18'd404: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=47;
   mapp<=64;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=12207;
 end   
18'd405: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=44;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd406: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd407: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=57;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd408: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd409: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd410: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd411: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd412: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd413: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11767;
 end   
18'd542: begin  
rid<=1;
end
18'd543: begin  
end
18'd544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd548: begin  
rid<=0;
end
18'd601: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=29;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1189;
 end   
18'd602: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd742: begin  
rid<=1;
end
18'd743: begin  
end
18'd744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd745: begin  
rid<=0;
end
18'd801: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=46;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11128;
 end   
18'd802: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=5;
   mapp<=90;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=17786;
 end   
18'd803: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=90;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd804: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=29;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd805: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=70;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd806: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=50;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd807: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=6;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd808: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=1;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd809: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd810: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd811: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd812: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd813: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11128;
 end   
18'd814: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11128;
 end   
18'd815: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11128;
 end   
18'd816: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11128;
 end   
18'd817: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11128;
 end   
18'd942: begin  
rid<=1;
end
18'd943: begin  
end
18'd944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd946: begin  
rid<=0;
end
18'd1001: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=76;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10707;
 end   
18'd1002: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=31;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd1003: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=8;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd1004: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=44;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd1005: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=39;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd1006: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=26;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd1007: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=23;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd1008: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd1009: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd1010: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd1011: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd1012: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd1013: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10707;
 end   
18'd1014: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10707;
 end   
18'd1142: begin  
rid<=1;
end
18'd1143: begin  
end
18'd1144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd1145: begin  
rid<=0;
end
18'd1201: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=15;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=270;
 end   
18'd1202: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=82;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=1240;
 end   
18'd1203: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=29;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=455;
 end   
18'd1204: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=41;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=645;
 end   
18'd1205: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=33;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=535;
 end   
18'd1206: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd1342: begin  
rid<=1;
end
18'd1343: begin  
end
18'd1344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd1345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd1346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd1347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd1348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd1349: begin  
rid<=0;
end
18'd1401: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=72;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4621;
 end   
18'd1402: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=70;
   mapp<=30;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7734;
 end   
18'd1403: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=29;
   mapp<=77;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8101;
 end   
18'd1404: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=6;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=8066;
 end   
18'd1405: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=73;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=11925;
 end   
18'd1406: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=86;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=9017;
 end   
18'd1407: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=21;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=5418;
 end   
18'd1408: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd1409: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd1410: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd1411: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd1412: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd1542: begin  
rid<=1;
end
18'd1543: begin  
end
18'd1544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd1545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd1546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd1547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd1548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd1549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd1550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd1551: begin  
rid<=0;
end
18'd1601: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=61;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=17109;
 end   
18'd1602: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=36;
   mapp<=12;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=14874;
 end   
18'd1603: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=55;
   mapp<=86;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=17549;
 end   
18'd1604: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=67;
   mapp<=90;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=16343;
 end   
18'd1605: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=55;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=13609;
 end   
18'd1606: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=74;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=16572;
 end   
18'd1607: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=31;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd1608: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=52;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd1609: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=50;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd1610: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd1611: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd1612: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd1613: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17109;
 end   
18'd1742: begin  
rid<=1;
end
18'd1743: begin  
end
18'd1744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd1745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd1746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd1747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd1748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd1749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd1750: begin  
rid<=0;
end
18'd1801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=57;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7110;
 end   
18'd1802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=87;
   mapp<=66;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6382;
 end   
18'd1803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=30;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=2339;
 end   
18'd1804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=7;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=8346;
 end   
18'd1805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=91;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=5836;
 end   
18'd1806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=7;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=3668;
 end   
18'd1807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd1808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd1809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd1942: begin  
rid<=1;
end
18'd1943: begin  
end
18'd1944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd1945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd1946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd1947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd1948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd1949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd1950: begin  
rid<=0;
end
18'd2001: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=9;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=405;
 end   
18'd2002: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=9;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=415;
 end   
18'd2003: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=58;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=2630;
 end   
18'd2004: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=21;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=975;
 end   
18'd2005: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=88;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=4000;
 end   
18'd2006: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=22;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=1040;
 end   
18'd2007: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=46;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=2130;
 end   
18'd2008: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=6;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=340;
 end   
18'd2009: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=30;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=1430;
 end   
18'd2010: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=13;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[9]<=675;
 end   
18'd2011: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=68;
   mapp<=0;
   pp<=100;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[10]<=3160;
 end   
18'd2012: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd2142: begin  
rid<=1;
end
18'd2143: begin  
end
18'd2144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd2145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd2146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd2147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd2148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd2149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd2150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd2151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd2152: begin  
check<=expctdoutput[8]-outcheck;
end
18'd2153: begin  
check<=expctdoutput[9]-outcheck;
end
18'd2154: begin  
check<=expctdoutput[10]-outcheck;
end
18'd2155: begin  
rid<=0;
end
18'd2201: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=2;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=23394;
 end   
18'd2202: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=50;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd2203: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=91;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd2204: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=36;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd2205: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=74;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd2206: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=20;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd2207: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=96;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd2208: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=21;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd2209: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=48;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd2210: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=99;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd2211: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd2212: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd2213: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23394;
 end   
18'd2214: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23394;
 end   
18'd2215: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23394;
 end   
18'd2216: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23394;
 end   
18'd2217: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23394;
 end   
18'd2218: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23394;
 end   
18'd2219: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23394;
 end   
18'd2220: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23394;
 end   
18'd2342: begin  
rid<=1;
end
18'd2343: begin  
end
18'd2344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd2345: begin  
rid<=0;
end
18'd2401: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=34;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2754;
 end   
18'd2402: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=53;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4303;
 end   
18'd2403: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=99;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8039;
 end   
18'd2404: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=18;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=1488;
 end   
18'd2405: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=38;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=3118;
 end   
18'd2406: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=50;
 end   
18'd2407: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=88;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=7188;
 end   
18'd2408: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=27;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=2257;
 end   
18'd2409: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=67;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=5507;
 end   
18'd2410: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=28;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[9]<=2358;
 end   
18'd2411: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd2542: begin  
rid<=1;
end
18'd2543: begin  
end
18'd2544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd2545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd2546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd2547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd2548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd2549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd2550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd2551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd2552: begin  
check<=expctdoutput[8]-outcheck;
end
18'd2553: begin  
check<=expctdoutput[9]-outcheck;
end
18'd2554: begin  
rid<=0;
end
18'd2601: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4119;
 end   
18'd2602: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=49;
   mapp<=7;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5381;
 end   
18'd2603: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=19;
   mapp<=21;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5868;
 end   
18'd2604: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=56;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd2605: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=98;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd2606: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=3;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd2607: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=24;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd2608: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=8;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd2609: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=44;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd2610: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd2611: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd2612: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd2613: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=4119;
 end   
18'd2614: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=4119;
 end   
18'd2615: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=4119;
 end   
18'd2616: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=4119;
 end   
18'd2617: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=4119;
 end   
18'd2618: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=4119;
 end   
18'd2619: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=4119;
 end   
18'd2620: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=4119;
 end   
18'd2742: begin  
rid<=1;
end
18'd2743: begin  
end
18'd2744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd2745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd2746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd2747: begin  
rid<=0;
end
18'd2801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=87;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7557;
 end   
18'd2802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=14;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7311;
 end   
18'd2803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=3;
   mapp<=85;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12594;
 end   
18'd2804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=48;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd2805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd2806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=58;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd2807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=18;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd2808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=80;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd2809: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd2810: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd2811: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd2812: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd2813: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7557;
 end   
18'd2814: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7557;
 end   
18'd2942: begin  
rid<=1;
end
18'd2943: begin  
end
18'd2944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd2945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd2946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd2947: begin  
rid<=0;
end
18'd3001: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=92;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=19386;
 end   
18'd3002: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=38;
   mapp<=89;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=17763;
 end   
18'd3003: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=79;
   mapp<=98;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=20361;
 end   
18'd3004: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=90;
   mapp<=9;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=10692;
 end   
18'd3005: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=57;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=13178;
 end   
18'd3006: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd3007: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd3008: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd3009: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd3010: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd3011: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd3012: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd3142: begin  
rid<=1;
end
18'd3143: begin  
end
18'd3144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd3145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd3146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd3147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd3148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd3149: begin  
rid<=0;
end
18'd3201: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=88;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8848;
 end   
18'd3202: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=56;
   mapp<=15;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5271;
 end   
18'd3203: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=11;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1051;
 end   
18'd3204: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=2;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=722;
 end   
18'd3205: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=34;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=4214;
 end   
18'd3206: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=72;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd3207: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd3208: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd3342: begin  
rid<=1;
end
18'd3343: begin  
end
18'd3344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd3345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd3346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd3347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd3348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd3349: begin  
rid<=0;
end
18'd3401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=75;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3450;
 end   
18'd3402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=62;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=4660;
 end   
18'd3403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=86;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=6470;
 end   
18'd3404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd3542: begin  
rid<=1;
end
18'd3543: begin  
end
18'd3544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd3545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd3546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd3547: begin  
rid<=0;
end
18'd3601: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=76;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15915;
 end   
18'd3602: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=92;
   mapp<=44;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=19649;
 end   
18'd3603: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=89;
   mapp<=16;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=19672;
 end   
18'd3604: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=75;
   mapp<=81;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=21237;
 end   
18'd3605: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=12;
   mapp<=98;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=16814;
 end   
18'd3606: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=22;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=16392;
 end   
18'd3607: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd3608: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd3609: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd3610: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd3611: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd3612: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd3613: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15915;
 end   
18'd3614: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15915;
 end   
18'd3615: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15915;
 end   
18'd3742: begin  
rid<=1;
end
18'd3743: begin  
end
18'd3744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd3745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd3746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd3747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd3748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd3749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd3750: begin  
rid<=0;
end
18'd3801: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=89;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5465;
 end   
18'd3802: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=55;
   mapp<=69;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11530;
 end   
18'd3803: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=23;
   mapp<=61;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=10312;
 end   
18'd3804: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd3805: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd3806: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd3807: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd3808: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd3942: begin  
rid<=1;
end
18'd3943: begin  
end
18'd3944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd3945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd3946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd3947: begin  
rid<=0;
end
18'd4001: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=54;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16021;
 end   
18'd4002: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=21;
   mapp<=85;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10054;
 end   
18'd4003: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=89;
   mapp<=88;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=11163;
 end   
18'd4004: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=76;
   mapp<=26;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=9296;
 end   
18'd4005: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=17;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=7435;
 end   
18'd4006: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=57;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=11892;
 end   
18'd4007: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd4008: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd4009: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd4010: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd4011: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd4012: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd4013: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16021;
 end   
18'd4142: begin  
rid<=1;
end
18'd4143: begin  
end
18'd4144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd4145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd4146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd4147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd4148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd4149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd4150: begin  
rid<=0;
end
18'd4201: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=55;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5910;
 end   
18'd4202: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=34;
   mapp<=25;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4363;
 end   
18'd4203: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=49;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5553;
 end   
18'd4204: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=41;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd4205: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd4206: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd4342: begin  
rid<=1;
end
18'd4343: begin  
end
18'd4344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd4345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd4346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd4347: begin  
rid<=0;
end
18'd4401: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=49;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=18659;
 end   
18'd4402: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=37;
   mapp<=18;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=23021;
 end   
18'd4403: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=66;
   mapp<=53;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=26642;
 end   
18'd4404: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=49;
   mapp<=39;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=23556;
 end   
18'd4405: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=93;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd4406: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=95;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd4407: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd4408: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd4409: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd4410: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd4411: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd4412: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd4413: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18659;
 end   
18'd4414: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18659;
 end   
18'd4415: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18659;
 end   
18'd4542: begin  
rid<=1;
end
18'd4543: begin  
end
18'd4544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd4545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd4546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd4547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd4548: begin  
rid<=0;
end
18'd4601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=71;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6106;
 end   
18'd4602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=365;
 end   
18'd4603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=88;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=6268;
 end   
18'd4604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=82;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=5852;
 end   
18'd4605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=55;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=3945;
 end   
18'd4606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=34;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=2464;
 end   
18'd4607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=14;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=1054;
 end   
18'd4608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=1;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=141;
 end   
18'd4609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=16;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=1216;
 end   
18'd4610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd4742: begin  
rid<=1;
end
18'd4743: begin  
end
18'd4744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd4745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd4746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd4747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd4748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd4749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd4750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd4751: begin  
check<=expctdoutput[7]-outcheck;
end
18'd4752: begin  
check<=expctdoutput[8]-outcheck;
end
18'd4753: begin  
rid<=0;
end
18'd4801: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=55;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=715;
 end   
18'd4802: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=85;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1115;
 end   
18'd4803: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=53;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=709;
 end   
18'd4804: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=12;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=186;
 end   
18'd4805: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=8;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=144;
 end   
18'd4806: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=32;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=466;
 end   
18'd4807: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=45;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=645;
 end   
18'd4808: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=13;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=239;
 end   
18'd4809: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=56;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=808;
 end   
18'd4810: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=21;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[9]<=363;
 end   
18'd4811: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd4942: begin  
rid<=1;
end
18'd4943: begin  
end
18'd4944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd4945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd4946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd4947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd4948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd4949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd4950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd4951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd4952: begin  
check<=expctdoutput[8]-outcheck;
end
18'd4953: begin  
check<=expctdoutput[9]-outcheck;
end
18'd4954: begin  
rid<=0;
end
18'd5001: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=81;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6642;
 end   
18'd5002: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=44;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3618;
 end   
18'd5003: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=96;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=7892;
 end   
18'd5004: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=22;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=1834;
 end   
18'd5005: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=29;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=2418;
 end   
18'd5006: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=61;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=5052;
 end   
18'd5007: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=35;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=2930;
 end   
18'd5008: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=50;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=4170;
 end   
18'd5009: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd5142: begin  
rid<=1;
end
18'd5143: begin  
end
18'd5144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd5145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd5146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd5147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd5148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd5149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd5150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd5151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd5152: begin  
rid<=0;
end
18'd5201: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=49;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14110;
 end   
18'd5202: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=86;
   mapp<=59;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=19442;
 end   
18'd5203: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=13;
   mapp<=92;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12215;
 end   
18'd5204: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=74;
   mapp<=39;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=14087;
 end   
18'd5205: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=22;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd5206: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=68;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd5207: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd5208: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd5209: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd5210: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd5211: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd5212: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd5213: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14110;
 end   
18'd5214: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14110;
 end   
18'd5215: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14110;
 end   
18'd5342: begin  
rid<=1;
end
18'd5343: begin  
end
18'd5344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd5345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd5346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd5347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd5348: begin  
rid<=0;
end
18'd5401: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=77;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3369;
 end   
18'd5402: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=14;
   mapp<=58;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4994;
 end   
18'd5403: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=14;
   mapp<=91;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6524;
 end   
18'd5404: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=24;
   mapp<=2;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=10475;
 end   
18'd5405: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=34;
   mapp<=25;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=11997;
 end   
18'd5406: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=74;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=11781;
 end   
18'd5407: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=72;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=9160;
 end   
18'd5408: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=59;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd5409: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=33;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd5410: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd5411: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=87;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd5412: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd5413: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=3369;
 end   
18'd5414: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=3369;
 end   
18'd5415: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=3369;
 end   
18'd5416: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=3369;
 end   
18'd5542: begin  
rid<=1;
end
18'd5543: begin  
end
18'd5544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd5545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd5546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd5547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd5548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd5549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd5550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd5551: begin  
rid<=0;
end
18'd5601: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=85;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15130;
 end   
18'd5602: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=2;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd5603: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=80;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd5604: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=13;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd5605: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=27;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd5606: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=2;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd5607: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd5608: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd5609: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd5610: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd5611: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd5612: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd5742: begin  
rid<=1;
end
18'd5743: begin  
end
18'd5744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd5745: begin  
rid<=0;
end
18'd5801: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=32;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3247;
 end   
18'd5802: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=5;
   mapp<=43;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3645;
 end   
18'd5803: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=93;
   mapp<=24;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=7599;
 end   
18'd5804: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=23;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=6799;
 end   
18'd5805: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=72;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=10182;
 end   
18'd5806: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=61;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=2686;
 end   
18'd5807: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd5808: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd5809: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd5810: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd5811: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd5942: begin  
rid<=1;
end
18'd5943: begin  
end
18'd5944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd5945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd5946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd5947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd5948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd5949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd5950: begin  
rid<=0;
end
18'd6001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=70;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=24351;
 end   
18'd6002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=35;
   mapp<=42;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=20739;
 end   
18'd6003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=33;
   mapp<=22;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=24823;
 end   
18'd6004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=11;
   mapp<=86;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=25003;
 end   
18'd6005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=60;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd6006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=96;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd6007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=67;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd6008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=85;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd6009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd6010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd6011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd6012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd6013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24351;
 end   
18'd6014: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24351;
 end   
18'd6015: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24351;
 end   
18'd6016: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24351;
 end   
18'd6017: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24351;
 end   
18'd6018: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24351;
 end   
18'd6019: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24351;
 end   
18'd6142: begin  
rid<=1;
end
18'd6143: begin  
end
18'd6144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd6145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd6146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd6147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd6148: begin  
rid<=0;
end
18'd6201: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=78;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=29103;
 end   
18'd6202: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=93;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=21311;
 end   
18'd6203: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=51;
   mapp<=24;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=20452;
 end   
18'd6204: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=84;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd6205: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=18;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd6206: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=64;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd6207: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=19;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd6208: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=52;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd6209: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd6210: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd6211: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd6212: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd6213: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29103;
 end   
18'd6214: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29103;
 end   
18'd6215: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29103;
 end   
18'd6216: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29103;
 end   
18'd6217: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29103;
 end   
18'd6218: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29103;
 end   
18'd6219: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29103;
 end   
18'd6220: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29103;
 end   
18'd6342: begin  
rid<=1;
end
18'd6343: begin  
end
18'd6344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd6345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd6346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd6347: begin  
rid<=0;
end
18'd6401: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=15;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5699;
 end   
18'd6402: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=76;
   mapp<=10;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8767;
 end   
18'd6403: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=27;
   mapp<=57;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8938;
 end   
18'd6404: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=43;
   mapp<=70;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=6006;
 end   
18'd6405: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=58;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=8441;
 end   
18'd6406: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=64;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd6407: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=9;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd6408: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=82;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd6409: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd6410: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd6411: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd6412: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd6542: begin  
rid<=1;
end
18'd6543: begin  
end
18'd6544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd6545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd6546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd6547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd6548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd6549: begin  
rid<=0;
end
18'd6601: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=27;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7229;
 end   
18'd6602: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=29;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6891;
 end   
18'd6603: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=28;
   mapp<=74;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5757;
 end   
18'd6604: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=23;
   mapp<=25;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=5269;
 end   
18'd6605: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=20;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=7097;
 end   
18'd6606: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=2;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=9100;
 end   
18'd6607: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd6608: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd6609: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=96;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd6610: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd6611: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd6612: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd6613: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7229;
 end   
18'd6742: begin  
rid<=1;
end
18'd6743: begin  
end
18'd6744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd6745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd6746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd6747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd6748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd6749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd6750: begin  
rid<=0;
end
18'd6801: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=71;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15408;
 end   
18'd6802: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=11;
   mapp<=25;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9059;
 end   
18'd6803: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=47;
   mapp<=64;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9370;
 end   
18'd6804: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=53;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd6805: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=20;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd6806: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=90;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd6807: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=24;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd6808: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd6809: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd6810: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd6811: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd6812: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd6813: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15408;
 end   
18'd6814: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15408;
 end   
18'd6815: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15408;
 end   
18'd6816: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15408;
 end   
18'd6942: begin  
rid<=1;
end
18'd6943: begin  
end
18'd6944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd6945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd6946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd6947: begin  
rid<=0;
end
18'd7001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=13;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10199;
 end   
18'd7002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=58;
   mapp<=51;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10541;
 end   
18'd7003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=78;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd7004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=65;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd7005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=7;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd7006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=77;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd7007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd7008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd7009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd7010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd7011: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd7142: begin  
rid<=1;
end
18'd7143: begin  
end
18'd7144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd7145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd7146: begin  
rid<=0;
end
18'd7201: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=60;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2511;
 end   
18'd7202: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=57;
   mapp<=3;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2305;
 end   
18'd7203: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=24;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1187;
 end   
18'd7204: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=77;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=3057;
 end   
18'd7205: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=8;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=391;
 end   
18'd7206: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=13;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=818;
 end   
18'd7207: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=87;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=3456;
 end   
18'd7208: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=1;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=259;
 end   
18'd7209: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=50;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=2210;
 end   
18'd7210: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=60;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[9]<=2514;
 end   
18'd7211: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=28;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd7212: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd7213: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=2511;
 end   
18'd7342: begin  
rid<=1;
end
18'd7343: begin  
end
18'd7344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd7345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd7346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd7347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd7348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd7349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd7350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd7351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd7352: begin  
check<=expctdoutput[8]-outcheck;
end
18'd7353: begin  
check<=expctdoutput[9]-outcheck;
end
18'd7354: begin  
rid<=0;
end
18'd7401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=4;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2036;
 end   
18'd7402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=35;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3217;
 end   
18'd7403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=56;
   mapp<=11;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=3730;
 end   
18'd7404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=72;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=2643;
 end   
18'd7405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=50;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd7406: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd7407: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd7408: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd7409: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd7542: begin  
rid<=1;
end
18'd7543: begin  
end
18'd7544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd7545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd7546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd7547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd7548: begin  
rid<=0;
end
18'd7601: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=22;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16804;
 end   
18'd7602: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=17;
   mapp<=26;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=19435;
 end   
18'd7603: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=12;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd7604: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=17;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd7605: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=96;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd7606: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=85;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd7607: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=41;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd7608: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=23;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd7609: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=29;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd7610: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd7611: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd7612: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd7613: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16804;
 end   
18'd7614: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16804;
 end   
18'd7615: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16804;
 end   
18'd7616: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16804;
 end   
18'd7617: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16804;
 end   
18'd7618: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16804;
 end   
18'd7619: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16804;
 end   
18'd7742: begin  
rid<=1;
end
18'd7743: begin  
end
18'd7744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd7745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd7746: begin  
rid<=0;
end
18'd7801: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=54;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3186;
 end   
18'd7802: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=1738;
 end   
18'd7803: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=96;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=5204;
 end   
18'd7804: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=55;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=3000;
 end   
18'd7805: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=53;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=2902;
 end   
18'd7806: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=62;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=3398;
 end   
18'd7807: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=84;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=4596;
 end   
18'd7808: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=34;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=1906;
 end   
18'd7809: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd7942: begin  
rid<=1;
end
18'd7943: begin  
end
18'd7944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd7945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd7946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd7947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd7948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd7949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd7950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd7951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd7952: begin  
rid<=0;
end
18'd8001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=23;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14378;
 end   
18'd8002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=42;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=12912;
 end   
18'd8003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=54;
   mapp<=63;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=17533;
 end   
18'd8004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=11;
   mapp<=7;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=16378;
 end   
18'd8005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=41;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd8006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=75;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd8007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=59;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd8008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=25;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd8009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd8010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd8011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd8012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd8013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14378;
 end   
18'd8014: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14378;
 end   
18'd8015: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14378;
 end   
18'd8016: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14378;
 end   
18'd8017: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14378;
 end   
18'd8018: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14378;
 end   
18'd8019: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14378;
 end   
18'd8142: begin  
rid<=1;
end
18'd8143: begin  
end
18'd8144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd8145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd8146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd8147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd8148: begin  
rid<=0;
end
18'd8201: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=37;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=19305;
 end   
18'd8202: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=34;
   mapp<=34;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=18641;
 end   
18'd8203: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=56;
   mapp<=5;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=26716;
 end   
18'd8204: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=93;
   mapp<=83;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=20285;
 end   
18'd8205: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=76;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd8206: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=5;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd8207: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=62;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd8208: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd8209: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd8210: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd8211: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd8212: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd8213: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19305;
 end   
18'd8214: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19305;
 end   
18'd8215: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19305;
 end   
18'd8216: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19305;
 end   
18'd8217: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19305;
 end   
18'd8342: begin  
rid<=1;
end
18'd8343: begin  
end
18'd8344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd8345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd8346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd8347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd8348: begin  
rid<=0;
end
18'd8401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=52;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=18084;
 end   
18'd8402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=43;
   mapp<=13;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=21031;
 end   
18'd8403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=96;
   mapp<=41;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=24393;
 end   
18'd8404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=73;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd8405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=40;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd8406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=13;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd8407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=75;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd8408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=72;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd8409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=18;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd8410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd8411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd8412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd8413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18084;
 end   
18'd8414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18084;
 end   
18'd8415: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18084;
 end   
18'd8416: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18084;
 end   
18'd8417: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18084;
 end   
18'd8418: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18084;
 end   
18'd8419: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18084;
 end   
18'd8420: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18084;
 end   
18'd8542: begin  
rid<=1;
end
18'd8543: begin  
end
18'd8544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd8545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd8546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd8547: begin  
rid<=0;
end
18'd8601: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=88;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=25438;
 end   
18'd8602: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=85;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd8603: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=90;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd8604: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=97;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd8605: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=89;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd8606: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=90;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd8607: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd8608: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd8609: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd8610: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd8611: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd8612: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd8742: begin  
rid<=1;
end
18'd8743: begin  
end
18'd8744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd8745: begin  
rid<=0;
end
18'd8801: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=81;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6211;
 end   
18'd8802: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=3;
   mapp<=51;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10167;
 end   
18'd8803: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=29;
   mapp<=40;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8171;
 end   
18'd8804: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=75;
   mapp<=44;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=9944;
 end   
18'd8805: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=8;
   mapp<=58;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=13494;
 end   
18'd8806: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=35;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=6617;
 end   
18'd8807: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd8808: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd8809: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd8810: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd8811: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd8812: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd8813: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6211;
 end   
18'd8814: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6211;
 end   
18'd8815: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6211;
 end   
18'd8942: begin  
rid<=1;
end
18'd8943: begin  
end
18'd8944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd8945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd8946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd8947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd8948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd8949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd8950: begin  
rid<=0;
end
18'd9001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=77;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9676;
 end   
18'd9002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=15;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7478;
 end   
18'd9003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=83;
   mapp<=61;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=10683;
 end   
18'd9004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=27;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=6517;
 end   
18'd9005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=67;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=8221;
 end   
18'd9006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=41;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=6962;
 end   
18'd9007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=29;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=3972;
 end   
18'd9008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=40;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=9487;
 end   
18'd9009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=13;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=2274;
 end   
18'd9010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd9011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd9012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd9013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9676;
 end   
18'd9014: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9676;
 end   
18'd9142: begin  
rid<=1;
end
18'd9143: begin  
end
18'd9144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd9145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd9146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd9147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd9148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd9149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd9150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd9151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd9152: begin  
check<=expctdoutput[8]-outcheck;
end
18'd9153: begin  
rid<=0;
end
18'd9201: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=75;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1886;
 end   
18'd9202: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=86;
   mapp<=1;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7997;
 end   
18'd9203: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=92;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=11994;
 end   
18'd9204: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=59;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=10475;
 end   
18'd9205: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=70;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=7698;
 end   
18'd9206: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=28;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=4472;
 end   
18'd9207: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=27;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=9309;
 end   
18'd9208: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd9209: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd9210: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd9342: begin  
rid<=1;
end
18'd9343: begin  
end
18'd9344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd9345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd9346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd9347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd9348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd9349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd9350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd9351: begin  
rid<=0;
end
18'd9401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=40;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3480;
 end   
18'd9402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=47;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=1890;
 end   
18'd9403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=4;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=180;
 end   
18'd9404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=3;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=150;
 end   
18'd9405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=21;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=880;
 end   
18'd9406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=63;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=2570;
 end   
18'd9407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=6;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=300;
 end   
18'd9408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=63;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=2590;
 end   
18'd9409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=10;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=480;
 end   
18'd9410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=71;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[9]<=2930;
 end   
18'd9411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=89;
   pp<=100;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[10]<=3660;
 end   
18'd9412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd9542: begin  
rid<=1;
end
18'd9543: begin  
end
18'd9544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd9545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd9546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd9547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd9548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd9549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd9550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd9551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd9552: begin  
check<=expctdoutput[8]-outcheck;
end
18'd9553: begin  
check<=expctdoutput[9]-outcheck;
end
18'd9554: begin  
check<=expctdoutput[10]-outcheck;
end
18'd9555: begin  
rid<=0;
end
18'd9601: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=3;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=57;
 end   
18'd9602: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=13;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=49;
 end   
18'd9603: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=91;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=293;
 end   
18'd9604: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=4;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=42;
 end   
18'd9605: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=18;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=94;
 end   
18'd9606: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=32;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=146;
 end   
18'd9607: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=50;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=210;
 end   
18'd9608: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=5;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=85;
 end   
18'd9609: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=75;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=305;
 end   
18'd9610: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=39;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[9]<=207;
 end   
18'd9611: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd9742: begin  
rid<=1;
end
18'd9743: begin  
end
18'd9744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd9745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd9746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd9747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd9748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd9749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd9750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd9751: begin  
check<=expctdoutput[7]-outcheck;
end
18'd9752: begin  
check<=expctdoutput[8]-outcheck;
end
18'd9753: begin  
check<=expctdoutput[9]-outcheck;
end
18'd9754: begin  
rid<=0;
end
18'd9801: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=13;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=611;
 end   
18'd9802: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=84;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=1102;
 end   
18'd9803: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=48;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=644;
 end   
18'd9804: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=71;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=953;
 end   
18'd9805: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=64;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=872;
 end   
18'd9806: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd9942: begin  
rid<=1;
end
18'd9943: begin  
end
18'd9944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd9945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd9946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd9947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd9948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd9949: begin  
rid<=0;
end
18'd10001: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=40;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13578;
 end   
18'd10002: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=45;
   mapp<=46;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11898;
 end   
18'd10003: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=8;
   mapp<=78;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=16214;
 end   
18'd10004: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=18;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd10005: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=70;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd10006: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=1;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd10007: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=23;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd10008: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=32;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd10009: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd10010: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd10011: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd10012: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd10013: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13578;
 end   
18'd10014: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13578;
 end   
18'd10015: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13578;
 end   
18'd10016: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13578;
 end   
18'd10017: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13578;
 end   
18'd10018: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13578;
 end   
18'd10142: begin  
rid<=1;
end
18'd10143: begin  
end
18'd10144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd10145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd10146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd10147: begin  
rid<=0;
end
18'd10201: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=15;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7803;
 end   
18'd10202: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=65;
   mapp<=70;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6393;
 end   
18'd10203: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=28;
   mapp<=63;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=3372;
 end   
18'd10204: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=43;
   mapp<=1;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=2045;
 end   
18'd10205: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=47;
   mapp<=3;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=5579;
 end   
18'd10206: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd10207: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd10208: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd10209: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd10210: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd10211: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd10212: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd10213: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7803;
 end   
18'd10214: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7803;
 end   
18'd10342: begin  
rid<=1;
end
18'd10343: begin  
end
18'd10344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd10345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd10346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd10347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd10348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd10349: begin  
rid<=0;
end
18'd10401: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=58;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=23838;
 end   
18'd10402: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=54;
   mapp<=9;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=22294;
 end   
18'd10403: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=88;
   mapp<=63;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=24248;
 end   
18'd10404: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=46;
   mapp<=49;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=21485;
 end   
18'd10405: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=90;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd10406: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=49;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd10407: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=43;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd10408: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd10409: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd10410: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd10411: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd10412: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd10413: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23838;
 end   
18'd10414: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23838;
 end   
18'd10415: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23838;
 end   
18'd10416: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23838;
 end   
18'd10417: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23838;
 end   
18'd10542: begin  
rid<=1;
end
18'd10543: begin  
end
18'd10544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd10545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd10546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd10547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd10548: begin  
rid<=0;
end
18'd10601: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=83;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6329;
 end   
18'd10602: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=35;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6831;
 end   
18'd10603: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd10604: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd10605: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd10742: begin  
rid<=1;
end
18'd10743: begin  
end
18'd10744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd10745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd10746: begin  
rid<=0;
end
18'd10801: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=66;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8368;
 end   
18'd10802: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=44;
   mapp<=53;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8215;
 end   
18'd10803: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=55;
   mapp<=29;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8205;
 end   
18'd10804: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=18;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd10805: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=26;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd10806: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=11;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd10807: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd10808: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd10809: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd10810: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd10811: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd10812: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd10813: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8368;
 end   
18'd10814: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8368;
 end   
18'd10942: begin  
rid<=1;
end
18'd10943: begin  
end
18'd10944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd10945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd10946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd10947: begin  
rid<=0;
end
18'd11001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=64;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11044;
 end   
18'd11002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=42;
   mapp<=49;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9943;
 end   
18'd11003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=75;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd11004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=13;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd11005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=42;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd11006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=96;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd11007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd11008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd11009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd11010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd11011: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd11142: begin  
rid<=1;
end
18'd11143: begin  
end
18'd11144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd11145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd11146: begin  
rid<=0;
end
18'd11201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=4;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2380;
 end   
18'd11202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=5;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd11203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=26;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd11204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=12;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd11205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd11206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd11207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd11208: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd11342: begin  
rid<=1;
end
18'd11343: begin  
end
18'd11344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd11345: begin  
rid<=0;
end
18'd11401: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=94;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12006;
 end   
18'd11402: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=56;
   mapp<=36;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9524;
 end   
18'd11403: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=52;
   mapp<=36;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=10196;
 end   
18'd11404: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=36;
   mapp<=41;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=9155;
 end   
18'd11405: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=38;
   mapp<=14;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=8491;
 end   
18'd11406: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=82;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd11407: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=55;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd11408: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=15;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd11409: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=31;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd11410: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd11411: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd11412: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd11413: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12006;
 end   
18'd11414: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12006;
 end   
18'd11542: begin  
rid<=1;
end
18'd11543: begin  
end
18'd11544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd11545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd11546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd11547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd11548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd11549: begin  
rid<=0;
end
18'd11601: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=90;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8018;
 end   
18'd11602: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=50;
   mapp<=11;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11198;
 end   
18'd11603: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=62;
   mapp<=37;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9943;
 end   
18'd11604: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=34;
   mapp<=86;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=5240;
 end   
18'd11605: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=93;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=8012;
 end   
18'd11606: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=53;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=4163;
 end   
18'd11607: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=16;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=6660;
 end   
18'd11608: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=52;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=6590;
 end   
18'd11609: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=8;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd11610: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd11611: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=33;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd11612: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd11613: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8018;
 end   
18'd11614: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8018;
 end   
18'd11615: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8018;
 end   
18'd11742: begin  
rid<=1;
end
18'd11743: begin  
end
18'd11744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd11745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd11746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd11747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd11748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd11749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd11750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd11751: begin  
check<=expctdoutput[7]-outcheck;
end
18'd11752: begin  
rid<=0;
end
18'd11801: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=80;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2774;
 end   
18'd11802: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=18;
   mapp<=3;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1258;
 end   
18'd11803: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=56;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=5364;
 end   
18'd11804: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=48;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=4302;
 end   
18'd11805: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=24;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=2266;
 end   
18'd11806: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=17;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=1644;
 end   
18'd11807: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=13;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=1262;
 end   
18'd11808: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=9;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=1294;
 end   
18'd11809: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=28;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=2320;
 end   
18'd11810: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd11811: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd11812: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd11942: begin  
rid<=1;
end
18'd11943: begin  
end
18'd11944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd11945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd11946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd11947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd11948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd11949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd11950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd11951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd11952: begin  
check<=expctdoutput[8]-outcheck;
end
18'd11953: begin  
rid<=0;
end
18'd12001: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=2;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15903;
 end   
18'd12002: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=61;
   mapp<=61;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11477;
 end   
18'd12003: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=89;
   mapp<=64;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9897;
 end   
18'd12004: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=48;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd12005: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=82;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd12006: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd12007: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd12008: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd12009: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd12010: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd12011: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd12012: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd12142: begin  
rid<=1;
end
18'd12143: begin  
end
18'd12144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd12145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd12146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd12147: begin  
rid<=0;
end
18'd12201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=31;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2552;
 end   
18'd12202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=69;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2903;
 end   
18'd12203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=78;
   mapp<=23;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1882;
 end   
18'd12204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=59;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=1663;
 end   
18'd12205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=8;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=1871;
 end   
18'd12206: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=19;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd12207: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=71;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd12208: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd12209: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd12210: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd12342: begin  
rid<=1;
end
18'd12343: begin  
end
18'd12344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd12345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd12346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd12347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd12348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd12349: begin  
rid<=0;
end
18'd12401: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=22;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1782;
 end   
18'd12402: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=4;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=98;
 end   
18'd12403: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=92;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=2044;
 end   
18'd12404: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=85;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=1900;
 end   
18'd12405: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=13;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=326;
 end   
18'd12406: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=98;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=2206;
 end   
18'd12407: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=89;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=2018;
 end   
18'd12408: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd12542: begin  
rid<=1;
end
18'd12543: begin  
end
18'd12544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd12545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd12546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd12547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd12548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd12549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd12550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd12551: begin  
rid<=0;
end
18'd12601: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=69;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11923;
 end   
18'd12602: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=58;
   mapp<=61;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=19899;
 end   
18'd12603: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=34;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=16296;
 end   
18'd12604: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=71;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd12605: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=64;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd12606: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=17;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd12607: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=15;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd12608: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=55;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd12609: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd12610: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd12611: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd12612: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd12613: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11923;
 end   
18'd12614: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11923;
 end   
18'd12615: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11923;
 end   
18'd12616: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11923;
 end   
18'd12617: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11923;
 end   
18'd12618: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11923;
 end   
18'd12742: begin  
rid<=1;
end
18'd12743: begin  
end
18'd12744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd12745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd12746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd12747: begin  
rid<=0;
end
18'd12801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=10;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15280;
 end   
18'd12802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=84;
   mapp<=12;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=19185;
 end   
18'd12803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=74;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd12804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=80;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd12805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=15;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd12806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd12807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd12808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd12809: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd12810: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd12811: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd12942: begin  
rid<=1;
end
18'd12943: begin  
end
18'd12944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd12945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd12946: begin  
rid<=0;
end
18'd13001: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=98;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8117;
 end   
18'd13002: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=73;
   mapp<=79;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8827;
 end   
18'd13003: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=88;
   mapp<=10;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=7743;
 end   
18'd13004: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=77;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=4273;
 end   
18'd13005: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=32;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=5834;
 end   
18'd13006: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=56;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=8051;
 end   
18'd13007: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd13008: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=13;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd13009: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd13010: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd13011: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd13142: begin  
rid<=1;
end
18'd13143: begin  
end
18'd13144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd13145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd13146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd13147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd13148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd13149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd13150: begin  
rid<=0;
end
18'd13201: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=71;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=26138;
 end   
18'd13202: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=33;
   mapp<=23;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=17460;
 end   
18'd13203: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=67;
   mapp<=63;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=20007;
 end   
18'd13204: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=53;
   mapp<=28;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=22541;
 end   
18'd13205: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=95;
   mapp<=84;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=25448;
 end   
18'd13206: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=68;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd13207: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd13208: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd13209: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd13210: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd13211: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd13212: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd13213: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26138;
 end   
18'd13214: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26138;
 end   
18'd13215: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26138;
 end   
18'd13216: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26138;
 end   
18'd13342: begin  
rid<=1;
end
18'd13343: begin  
end
18'd13344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd13345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd13346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd13347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd13348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd13349: begin  
rid<=0;
end
18'd13401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=9;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13339;
 end   
18'd13402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=93;
   mapp<=50;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=14847;
 end   
18'd13403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=86;
   mapp<=98;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8082;
 end   
18'd13404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=80;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=7952;
 end   
18'd13405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=16;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=9520;
 end   
18'd13406: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=49;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=7565;
 end   
18'd13407: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=67;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd13408: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=28;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd13409: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd13410: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd13411: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd13542: begin  
rid<=1;
end
18'd13543: begin  
end
18'd13544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd13545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd13546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd13547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd13548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd13549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd13550: begin  
rid<=0;
end
18'd13601: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=26;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5458;
 end   
18'd13602: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=66;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5601;
 end   
18'd13603: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=87;
   mapp<=26;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5932;
 end   
18'd13604: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=81;
   mapp<=16;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=4803;
 end   
18'd13605: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=64;
   mapp<=16;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=5148;
 end   
18'd13606: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=40;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=3194;
 end   
18'd13607: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=86;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=4943;
 end   
18'd13608: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=21;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd13609: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd13610: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=21;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd13611: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=64;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd13612: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd13613: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5458;
 end   
18'd13614: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5458;
 end   
18'd13615: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5458;
 end   
18'd13616: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5458;
 end   
18'd13742: begin  
rid<=1;
end
18'd13743: begin  
end
18'd13744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd13745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd13746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd13747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd13748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd13749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd13750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd13751: begin  
rid<=0;
end
18'd13801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=23;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6175;
 end   
18'd13802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=31;
   mapp<=73;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3404;
 end   
18'd13803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=6;
   mapp<=24;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6259;
 end   
18'd13804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=68;
   mapp<=41;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=7152;
 end   
18'd13805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=18;
   mapp<=45;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=5066;
 end   
18'd13806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=2;
   mapp<=62;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=6826;
 end   
18'd13807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=7;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd13808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=7;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd13809: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=81;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd13810: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd13811: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=36;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd13812: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd13813: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6175;
 end   
18'd13814: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6175;
 end   
18'd13815: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6175;
 end   
18'd13816: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6175;
 end   
18'd13817: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6175;
 end   
18'd13942: begin  
rid<=1;
end
18'd13943: begin  
end
18'd13944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd13945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd13946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd13947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd13948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd13949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd13950: begin  
rid<=0;
end
18'd14001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=91;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3563;
 end   
18'd14002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=12;
   mapp<=84;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11116;
 end   
18'd14003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=31;
   mapp<=56;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9079;
 end   
18'd14004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=90;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=12312;
 end   
18'd14005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=93;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=11267;
 end   
18'd14006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=96;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=11084;
 end   
18'd14007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=52;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=6835;
 end   
18'd14008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=54;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=5772;
 end   
18'd14009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=45;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=5759;
 end   
18'd14010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd14011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd14012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd14013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=3563;
 end   
18'd14014: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=3563;
 end   
18'd14142: begin  
rid<=1;
end
18'd14143: begin  
end
18'd14144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd14145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd14146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd14147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd14148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd14149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd14150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd14151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd14152: begin  
check<=expctdoutput[8]-outcheck;
end
18'd14153: begin  
rid<=0;
end
18'd14201: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=23;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=18629;
 end   
18'd14202: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=18;
   mapp<=22;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=23482;
 end   
18'd14203: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=66;
   mapp<=4;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=20335;
 end   
18'd14204: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=59;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd14205: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=98;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd14206: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=86;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd14207: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd14208: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd14209: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd14210: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd14211: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd14212: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd14213: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18629;
 end   
18'd14214: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18629;
 end   
18'd14342: begin  
rid<=1;
end
18'd14343: begin  
end
18'd14344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd14345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd14346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd14347: begin  
rid<=0;
end
18'd14401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=98;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14174;
 end   
18'd14402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=30;
   mapp<=58;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13472;
 end   
18'd14403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=92;
   mapp<=22;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=13970;
 end   
18'd14404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=46;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=14368;
 end   
18'd14405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=78;
   mapp<=92;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=16990;
 end   
18'd14406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=37;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=8906;
 end   
18'd14407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=25;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=9802;
 end   
18'd14408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd14409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd14410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd14411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd14412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd14413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14174;
 end   
18'd14414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14174;
 end   
18'd14415: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14174;
 end   
18'd14416: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14174;
 end   
18'd14542: begin  
rid<=1;
end
18'd14543: begin  
end
18'd14544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd14545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd14546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd14547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd14548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd14549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd14550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd14551: begin  
rid<=0;
end
18'd14601: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=97;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11482;
 end   
18'd14602: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=28;
   mapp<=82;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=12909;
 end   
18'd14603: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=51;
   mapp<=40;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=11147;
 end   
18'd14604: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=16;
   mapp<=15;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=8899;
 end   
18'd14605: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=30;
   mapp<=75;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=15954;
 end   
18'd14606: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=62;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=11868;
 end   
18'd14607: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd14608: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd14609: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd14610: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd14611: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd14612: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd14613: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11482;
 end   
18'd14614: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11482;
 end   
18'd14615: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11482;
 end   
18'd14742: begin  
rid<=1;
end
18'd14743: begin  
end
18'd14744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd14745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd14746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd14747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd14748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd14749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd14750: begin  
rid<=0;
end
18'd14801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=62;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16569;
 end   
18'd14802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=55;
   mapp<=29;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=17501;
 end   
18'd14803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=75;
   mapp<=20;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=18460;
 end   
18'd14804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=92;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd14805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=61;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd14806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=54;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd14807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=98;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd14808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=46;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd14809: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd14810: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd14811: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd14812: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd14813: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16569;
 end   
18'd14814: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16569;
 end   
18'd14942: begin  
rid<=1;
end
18'd14943: begin  
end
18'd14944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd14945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd14946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd14947: begin  
rid<=0;
end
18'd15001: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=63;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11289;
 end   
18'd15002: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=75;
   mapp<=69;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8443;
 end   
18'd15003: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=15;
   mapp<=38;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5639;
 end   
18'd15004: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=21;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=7623;
 end   
18'd15005: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=75;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=8739;
 end   
18'd15006: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=15;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=4594;
 end   
18'd15007: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=28;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd15008: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd15009: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd15010: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd15011: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd15142: begin  
rid<=1;
end
18'd15143: begin  
end
18'd15144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd15145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd15146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd15147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd15148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd15149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd15150: begin  
rid<=0;
end
18'd15201: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=50;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7241;
 end   
18'd15202: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=33;
   mapp<=57;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6671;
 end   
18'd15203: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=25;
   mapp<=62;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6223;
 end   
18'd15204: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=10;
   mapp<=61;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=5787;
 end   
18'd15205: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=24;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=4882;
 end   
18'd15206: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=49;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=5757;
 end   
18'd15207: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd15208: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd15209: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd15210: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd15211: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd15212: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd15213: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7241;
 end   
18'd15342: begin  
rid<=1;
end
18'd15343: begin  
end
18'd15344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd15345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd15346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd15347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd15348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd15349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd15350: begin  
rid<=0;
end
18'd15401: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=14;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5510;
 end   
18'd15402: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=64;
   mapp<=78;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7054;
 end   
18'd15403: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=93;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=3626;
 end   
18'd15404: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd15405: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd15406: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd15542: begin  
rid<=1;
end
18'd15543: begin  
end
18'd15544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd15545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd15546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd15547: begin  
rid<=0;
end
18'd15601: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=85;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13034;
 end   
18'd15602: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=52;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13421;
 end   
18'd15603: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=73;
   mapp<=37;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=18814;
 end   
18'd15604: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=52;
   mapp<=4;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=16257;
 end   
18'd15605: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=94;
   mapp<=37;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=20719;
 end   
18'd15606: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=76;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd15607: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=26;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd15608: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd15609: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd15610: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd15611: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd15612: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd15613: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13034;
 end   
18'd15614: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13034;
 end   
18'd15615: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13034;
 end   
18'd15616: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13034;
 end   
18'd15617: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13034;
 end   
18'd15618: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13034;
 end   
18'd15742: begin  
rid<=1;
end
18'd15743: begin  
end
18'd15744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd15745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd15746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd15747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd15748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd15749: begin  
rid<=0;
end
18'd15801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=41;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8425;
 end   
18'd15802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=89;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11447;
 end   
18'd15803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=19;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd15804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=65;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd15805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=5;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd15806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd15807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd15808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd15809: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd15810: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd15811: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd15942: begin  
rid<=1;
end
18'd15943: begin  
end
18'd15944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd15945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd15946: begin  
rid<=0;
end
18'd16001: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=9;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1305;
 end   
18'd16002: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=15;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6225;
 end   
18'd16003: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=95;
   mapp<=9;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6371;
 end   
18'd16004: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=64;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=9441;
 end   
18'd16005: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=66;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=7664;
 end   
18'd16006: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd16007: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd16008: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd16009: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd16010: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd16142: begin  
rid<=1;
end
18'd16143: begin  
end
18'd16144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd16145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd16146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd16147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd16148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd16149: begin  
rid<=0;
end
18'd16201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=31;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8555;
 end   
18'd16202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=68;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8374;
 end   
18'd16203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=26;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd16204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd16205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd16206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd16207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd16342: begin  
rid<=1;
end
18'd16343: begin  
end
18'd16344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd16345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd16346: begin  
rid<=0;
end
18'd16401: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=2;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16756;
 end   
18'd16402: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=55;
   mapp<=79;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=18453;
 end   
18'd16403: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=60;
   mapp<=10;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=22738;
 end   
18'd16404: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=74;
   mapp<=52;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=23296;
 end   
18'd16405: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=72;
   mapp<=82;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=22317;
 end   
18'd16406: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=21;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd16407: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd16408: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd16409: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd16410: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd16411: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd16412: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd16413: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16756;
 end   
18'd16414: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16756;
 end   
18'd16415: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16756;
 end   
18'd16416: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16756;
 end   
18'd16542: begin  
rid<=1;
end
18'd16543: begin  
end
18'd16544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd16545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd16546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd16547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd16548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd16549: begin  
rid<=0;
end
18'd16601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=12;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14415;
 end   
18'd16602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=72;
   mapp<=89;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11041;
 end   
18'd16603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=39;
   mapp<=5;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=15850;
 end   
18'd16604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=28;
   mapp<=95;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=16762;
 end   
18'd16605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=12;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd16606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=62;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd16607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd16608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd16609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd16610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd16611: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd16612: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd16613: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14415;
 end   
18'd16614: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14415;
 end   
18'd16615: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14415;
 end   
18'd16742: begin  
rid<=1;
end
18'd16743: begin  
end
18'd16744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd16745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd16746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd16747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd16748: begin  
rid<=0;
end
18'd16801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=86;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5899;
 end   
18'd16802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=19;
   mapp<=8;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4392;
 end   
18'd16803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=58;
   mapp<=23;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5550;
 end   
18'd16804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=45;
   mapp<=59;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=4917;
 end   
18'd16805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=6;
   mapp<=34;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=8087;
 end   
18'd16806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=66;
   mapp<=4;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=11095;
 end   
18'd16807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd16808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=67;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd16809: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=92;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd16810: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=87;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd16811: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=32;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd16812: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd16813: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5899;
 end   
18'd16814: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5899;
 end   
18'd16815: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5899;
 end   
18'd16816: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5899;
 end   
18'd16817: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5899;
 end   
18'd16942: begin  
rid<=1;
end
18'd16943: begin  
end
18'd16944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd16945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd16946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd16947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd16948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd16949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd16950: begin  
rid<=0;
end
18'd17001: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=18;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=27416;
 end   
18'd17002: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=76;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd17003: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=20;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd17004: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=11;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd17005: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=82;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd17006: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=56;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd17007: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=90;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd17008: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=25;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd17009: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=24;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd17010: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=86;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd17011: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd17012: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd17013: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=27416;
 end   
18'd17014: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=27416;
 end   
18'd17015: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=27416;
 end   
18'd17016: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=27416;
 end   
18'd17017: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=27416;
 end   
18'd17018: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=27416;
 end   
18'd17019: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=27416;
 end   
18'd17020: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=27416;
 end   
18'd17142: begin  
rid<=1;
end
18'd17143: begin  
end
18'd17144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd17145: begin  
rid<=0;
end
18'd17201: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=26;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=19205;
 end   
18'd17202: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=71;
   mapp<=34;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=18778;
 end   
18'd17203: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=97;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd17204: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=12;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd17205: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=3;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd17206: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=27;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd17207: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=8;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd17208: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=45;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd17209: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=8;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd17210: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd17211: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd17212: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd17213: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19205;
 end   
18'd17214: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19205;
 end   
18'd17215: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19205;
 end   
18'd17216: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19205;
 end   
18'd17217: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19205;
 end   
18'd17218: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19205;
 end   
18'd17219: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19205;
 end   
18'd17342: begin  
rid<=1;
end
18'd17343: begin  
end
18'd17344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd17345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd17346: begin  
rid<=0;
end
18'd17401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=1;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2551;
 end   
18'd17402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=50;
   mapp<=43;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3207;
 end   
18'd17403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=28;
   mapp<=13;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=2179;
 end   
18'd17404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=11;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=3224;
 end   
18'd17405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=50;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=5193;
 end   
18'd17406: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=49;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=6521;
 end   
18'd17407: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=92;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=6683;
 end   
18'd17408: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=54;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=6088;
 end   
18'd17409: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=69;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=6961;
 end   
18'd17410: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=81;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd17411: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=65;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd17412: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd17413: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=2551;
 end   
18'd17414: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=2551;
 end   
18'd17542: begin  
rid<=1;
end
18'd17543: begin  
end
18'd17544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd17545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd17546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd17547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd17548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd17549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd17550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd17551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd17552: begin  
check<=expctdoutput[8]-outcheck;
end
18'd17553: begin  
rid<=0;
end
18'd17601: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=42;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=17108;
 end   
18'd17602: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=77;
   mapp<=34;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=14626;
 end   
18'd17603: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=77;
   mapp<=72;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=10968;
 end   
18'd17604: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=70;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd17605: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd17606: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd17607: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd17608: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd17609: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd17610: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd17742: begin  
rid<=1;
end
18'd17743: begin  
end
18'd17744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd17745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd17746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd17747: begin  
rid<=0;
end
18'd17801: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=10;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=26308;
 end   
18'd17802: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=82;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd17803: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=58;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd17804: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=26;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd17805: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=87;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd17806: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=70;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd17807: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=28;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd17808: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=51;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd17809: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=58;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd17810: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=13;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd17811: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd17812: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd17813: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26308;
 end   
18'd17814: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26308;
 end   
18'd17815: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26308;
 end   
18'd17816: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26308;
 end   
18'd17817: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26308;
 end   
18'd17818: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26308;
 end   
18'd17819: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26308;
 end   
18'd17820: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26308;
 end   
18'd17942: begin  
rid<=1;
end
18'd17943: begin  
end
18'd17944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd17945: begin  
rid<=0;
end
18'd18001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=34;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6918;
 end   
18'd18002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=41;
   mapp<=42;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10966;
 end   
18'd18003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=18;
   mapp<=10;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8108;
 end   
18'd18004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=3;
   mapp<=72;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=8756;
 end   
18'd18005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=67;
   mapp<=28;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=16340;
 end   
18'd18006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=65;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=13550;
 end   
18'd18007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=38;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=11292;
 end   
18'd18008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=81;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd18009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=57;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd18010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=50;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd18011: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=14;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd18012: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd18013: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6918;
 end   
18'd18014: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6918;
 end   
18'd18015: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6918;
 end   
18'd18016: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6918;
 end   
18'd18142: begin  
rid<=1;
end
18'd18143: begin  
end
18'd18144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd18145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd18146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd18147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd18148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd18149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd18150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd18151: begin  
rid<=0;
end
18'd18201: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=86;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10664;
 end   
18'd18202: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=86;
   mapp<=63;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10244;
 end   
18'd18203: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=56;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=5438;
 end   
18'd18204: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=7;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=7340;
 end   
18'd18205: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=78;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=14402;
 end   
18'd18206: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=89;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=10714;
 end   
18'd18207: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=35;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=8660;
 end   
18'd18208: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=65;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=12110;
 end   
18'd18209: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd18210: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd18211: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd18342: begin  
rid<=1;
end
18'd18343: begin  
end
18'd18344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd18345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd18346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd18347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd18348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd18349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd18350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd18351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd18352: begin  
rid<=0;
end
18'd18401: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=28;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=840;
 end   
18'd18402: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=0;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=1354;
 end   
18'd18403: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd18542: begin  
rid<=1;
end
18'd18543: begin  
end
18'd18544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd18545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd18546: begin  
rid<=0;
end
18'd18601: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=35;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2060;
 end   
18'd18602: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=10;
   mapp<=66;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6944;
 end   
18'd18603: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=99;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6422;
 end   
18'd18604: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd18605: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd18606: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd18742: begin  
rid<=1;
end
18'd18743: begin  
end
18'd18744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd18745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd18746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd18747: begin  
rid<=0;
end
18'd18801: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=44;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6672;
 end   
18'd18802: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=94;
   mapp<=52;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6646;
 end   
18'd18803: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=8;
   mapp<=69;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6191;
 end   
18'd18804: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=52;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=6138;
 end   
18'd18805: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=47;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd18806: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=32;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd18807: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd18808: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd18809: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd18942: begin  
rid<=1;
end
18'd18943: begin  
end
18'd18944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd18945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd18946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd18947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd18948: begin  
rid<=0;
end
18'd19001: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=23;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11218;
 end   
18'd19002: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=51;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8555;
 end   
18'd19003: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=74;
   mapp<=43;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5971;
 end   
18'd19004: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=33;
   mapp<=49;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=7893;
 end   
18'd19005: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=15;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=9062;
 end   
18'd19006: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=41;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=5928;
 end   
18'd19007: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=89;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=4579;
 end   
18'd19008: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd19009: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd19010: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd19011: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd19012: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd19013: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11218;
 end   
18'd19014: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11218;
 end   
18'd19142: begin  
rid<=1;
end
18'd19143: begin  
end
18'd19144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd19145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd19146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd19147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd19148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd19149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd19150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd19151: begin  
rid<=0;
end
18'd19201: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=78;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=18990;
 end   
18'd19202: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=31;
   mapp<=90;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=19097;
 end   
18'd19203: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=44;
   mapp<=97;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=18316;
 end   
18'd19204: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=40;
   mapp<=19;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=26738;
 end   
18'd19205: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=87;
   mapp<=80;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=20690;
 end   
18'd19206: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=99;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd19207: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=25;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd19208: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=83;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd19209: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd19210: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd19211: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd19212: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd19213: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18990;
 end   
18'd19214: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18990;
 end   
18'd19342: begin  
rid<=1;
end
18'd19343: begin  
end
18'd19344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd19345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd19346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd19347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd19348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd19349: begin  
rid<=0;
end
18'd19401: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=60;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3120;
 end   
18'd19402: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=0;
   mapp<=11;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=670;
 end   
18'd19403: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd19542: begin  
rid<=1;
end
18'd19543: begin  
end
18'd19544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd19545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd19546: begin  
rid<=0;
end
18'd19601: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=92;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14315;
 end   
18'd19602: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=10;
   mapp<=85;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10470;
 end   
18'd19603: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=49;
   mapp<=29;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=10431;
 end   
18'd19604: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=78;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd19605: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd19606: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd19607: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd19608: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd19609: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd19610: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd19742: begin  
rid<=1;
end
18'd19743: begin  
end
18'd19744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd19745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd19746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd19747: begin  
rid<=0;
end
18'd19801: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=82;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=31746;
 end   
18'd19802: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=78;
   mapp<=73;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=27384;
 end   
18'd19803: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=59;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd19804: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=18;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd19805: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=89;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd19806: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=59;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd19807: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=49;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd19808: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd19809: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd19810: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd19811: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd19812: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd19813: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=31746;
 end   
18'd19814: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=31746;
 end   
18'd19815: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=31746;
 end   
18'd19942: begin  
rid<=1;
end
18'd19943: begin  
end
18'd19944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd19945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd19946: begin  
rid<=0;
end
18'd20001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=11;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=21680;
 end   
18'd20002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=19;
   mapp<=8;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=15336;
 end   
18'd20003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=61;
   mapp<=67;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=22371;
 end   
18'd20004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=56;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd20005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=90;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd20006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=63;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd20007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=83;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd20008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=16;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd20009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=32;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd20010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd20011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd20012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd20013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21680;
 end   
18'd20014: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21680;
 end   
18'd20015: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21680;
 end   
18'd20016: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21680;
 end   
18'd20017: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21680;
 end   
18'd20018: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21680;
 end   
18'd20019: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21680;
 end   
18'd20020: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21680;
 end   
18'd20142: begin  
rid<=1;
end
18'd20143: begin  
end
18'd20144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd20145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd20146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd20147: begin  
rid<=0;
end
18'd20201: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=98;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11102;
 end   
18'd20202: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=32;
   mapp<=13;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11620;
 end   
18'd20203: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=87;
   mapp<=62;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=14388;
 end   
18'd20204: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=96;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=12663;
 end   
18'd20205: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=60;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=6748;
 end   
18'd20206: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=15;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=10261;
 end   
18'd20207: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=4;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=6752;
 end   
18'd20208: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=99;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=17884;
 end   
18'd20209: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd20210: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd20211: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd20212: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd20213: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11102;
 end   
18'd20342: begin  
rid<=1;
end
18'd20343: begin  
end
18'd20344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd20345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd20346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd20347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd20348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd20349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd20350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd20351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd20352: begin  
rid<=0;
end
18'd20401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=41;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4619;
 end   
18'd20402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=82;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd20403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=49;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd20404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd20405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd20406: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd20542: begin  
rid<=1;
end
18'd20543: begin  
end
18'd20544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd20545: begin  
rid<=0;
end
18'd20601: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=16;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1718;
 end   
18'd20602: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=78;
   mapp<=21;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7756;
 end   
18'd20603: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=95;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=9028;
 end   
18'd20604: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd20605: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd20606: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd20742: begin  
rid<=1;
end
18'd20743: begin  
end
18'd20744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd20745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd20746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd20747: begin  
rid<=0;
end
18'd20801: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=29;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13215;
 end   
18'd20802: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=81;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=16455;
 end   
18'd20803: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=95;
   mapp<=50;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=15707;
 end   
18'd20804: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=78;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd20805: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=76;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd20806: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=53;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd20807: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd20808: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd20809: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd20810: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd20942: begin  
rid<=1;
end
18'd20943: begin  
end
18'd20944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd20945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd20946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd20947: begin  
rid<=0;
end
18'd21001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=22;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12494;
 end   
18'd21002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=48;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9810;
 end   
18'd21003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=51;
   mapp<=8;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8339;
 end   
18'd21004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=86;
   mapp<=72;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=6361;
 end   
18'd21005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=43;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=8940;
 end   
18'd21006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=29;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=9558;
 end   
18'd21007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=14;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=14263;
 end   
18'd21008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=68;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=15125;
 end   
18'd21009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd21010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd21011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd21012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd21013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12494;
 end   
18'd21014: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12494;
 end   
18'd21015: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12494;
 end   
18'd21142: begin  
rid<=1;
end
18'd21143: begin  
end
18'd21144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd21145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd21146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd21147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd21148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd21149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd21150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd21151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd21152: begin  
rid<=0;
end
18'd21201: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=15;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1988;
 end   
18'd21202: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=49;
   mapp<=17;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1686;
 end   
18'd21203: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=29;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=1239;
 end   
18'd21204: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=16;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=3896;
 end   
18'd21205: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=74;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=5609;
 end   
18'd21206: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=91;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=4796;
 end   
18'd21207: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=69;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=1683;
 end   
18'd21208: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=12;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=2504;
 end   
18'd21209: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=46;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=5327;
 end   
18'd21210: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=93;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[9]<=5944;
 end   
18'd21211: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd21212: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd21213: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=1988;
 end   
18'd21342: begin  
rid<=1;
end
18'd21343: begin  
end
18'd21344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd21345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd21346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd21347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd21348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd21349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd21350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd21351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd21352: begin  
check<=expctdoutput[8]-outcheck;
end
18'd21353: begin  
check<=expctdoutput[9]-outcheck;
end
18'd21354: begin  
rid<=0;
end
18'd21401: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=83;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=21909;
 end   
18'd21402: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=94;
   mapp<=36;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=21304;
 end   
18'd21403: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=80;
   mapp<=51;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=24100;
 end   
18'd21404: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=97;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd21405: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=65;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd21406: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd21407: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd21408: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd21409: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd21410: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd21411: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd21412: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd21542: begin  
rid<=1;
end
18'd21543: begin  
end
18'd21544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd21545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd21546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd21547: begin  
rid<=0;
end
18'd21601: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=47;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=21797;
 end   
18'd21602: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=45;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd21603: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=70;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd21604: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=75;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd21605: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=89;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd21606: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=50;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd21607: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd21608: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd21609: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd21610: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd21611: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd21612: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd21742: begin  
rid<=1;
end
18'd21743: begin  
end
18'd21744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd21745: begin  
rid<=0;
end
18'd21801: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=14;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=910;
 end   
18'd21802: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd21942: begin  
rid<=1;
end
18'd21943: begin  
end
18'd21944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd21945: begin  
rid<=0;
end
18'd22001: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=67;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4256;
 end   
18'd22002: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=22;
   mapp<=96;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8586;
 end   
18'd22003: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=82;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd22004: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd22005: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd22142: begin  
rid<=1;
end
18'd22143: begin  
end
18'd22144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd22145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd22146: begin  
rid<=0;
end
18'd22201: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=76;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=18559;
 end   
18'd22202: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=59;
   mapp<=87;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=24757;
 end   
18'd22203: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=89;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd22204: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=22;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd22205: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=66;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd22206: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=86;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd22207: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=55;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd22208: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=28;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd22209: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=14;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd22210: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd22211: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd22212: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd22213: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18559;
 end   
18'd22214: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18559;
 end   
18'd22215: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18559;
 end   
18'd22216: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18559;
 end   
18'd22217: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18559;
 end   
18'd22218: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18559;
 end   
18'd22219: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18559;
 end   
18'd22342: begin  
rid<=1;
end
18'd22343: begin  
end
18'd22344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd22345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd22346: begin  
rid<=0;
end
18'd22401: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=21;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9454;
 end   
18'd22402: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=96;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11408;
 end   
18'd22403: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=81;
   mapp<=3;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=13197;
 end   
18'd22404: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=21;
   mapp<=61;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=17419;
 end   
18'd22405: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=55;
   mapp<=31;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=15385;
 end   
18'd22406: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=82;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=17895;
 end   
18'd22407: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd22408: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd22409: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd22410: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd22411: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd22412: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd22413: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9454;
 end   
18'd22414: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9454;
 end   
18'd22415: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9454;
 end   
18'd22542: begin  
rid<=1;
end
18'd22543: begin  
end
18'd22544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd22545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd22546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd22547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd22548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd22549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd22550: begin  
rid<=0;
end
18'd22601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=35;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=28253;
 end   
18'd22602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=43;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=28031;
 end   
18'd22603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=88;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd22604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=53;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd22605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=32;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd22606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=47;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd22607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=80;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd22608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=26;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd22609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=78;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd22610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=50;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd22611: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd22612: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd22613: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28253;
 end   
18'd22614: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28253;
 end   
18'd22615: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28253;
 end   
18'd22616: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28253;
 end   
18'd22617: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28253;
 end   
18'd22618: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28253;
 end   
18'd22619: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28253;
 end   
18'd22742: begin  
rid<=1;
end
18'd22743: begin  
end
18'd22744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd22745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd22746: begin  
rid<=0;
end
18'd22801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=73;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14447;
 end   
18'd22802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=74;
   mapp<=55;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9487;
 end   
18'd22803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=50;
   mapp<=63;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9453;
 end   
18'd22804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=16;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=9650;
 end   
18'd22805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=73;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=12133;
 end   
18'd22806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd22807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd22808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd22809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd22810: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd22942: begin  
rid<=1;
end
18'd22943: begin  
end
18'd22944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd22945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd22946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd22947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd22948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd22949: begin  
rid<=0;
end
18'd23001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=47;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=18604;
 end   
18'd23002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=90;
   mapp<=99;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=14125;
 end   
18'd23003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=71;
   mapp<=10;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=11423;
 end   
18'd23004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=5;
   mapp<=43;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=18990;
 end   
18'd23005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=72;
   mapp<=65;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=12903;
 end   
18'd23006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=72;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=17327;
 end   
18'd23007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=29;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=15777;
 end   
18'd23008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd23009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd23010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd23011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd23012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd23013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18604;
 end   
18'd23014: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18604;
 end   
18'd23015: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18604;
 end   
18'd23016: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18604;
 end   
18'd23142: begin  
rid<=1;
end
18'd23143: begin  
end
18'd23144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd23145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd23146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd23147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd23148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd23149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd23150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd23151: begin  
rid<=0;
end
18'd23201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=58;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7391;
 end   
18'd23202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=93;
   mapp<=65;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4678;
 end   
18'd23203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=6;
   mapp<=31;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6698;
 end   
18'd23204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=78;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=4896;
 end   
18'd23205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=48;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=3591;
 end   
18'd23206: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=6;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=6831;
 end   
18'd23207: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=71;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd23208: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=66;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd23209: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd23210: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd23211: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd23342: begin  
rid<=1;
end
18'd23343: begin  
end
18'd23344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd23345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd23346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd23347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd23348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd23349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd23350: begin  
rid<=0;
end
18'd23401: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=15;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=23197;
 end   
18'd23402: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=26;
   mapp<=94;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=29271;
 end   
18'd23403: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=84;
   mapp<=29;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=28492;
 end   
18'd23404: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=68;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd23405: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=6;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd23406: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=28;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd23407: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=97;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd23408: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=18;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd23409: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=90;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd23410: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=99;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd23411: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=85;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd23412: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd23413: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23197;
 end   
18'd23414: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23197;
 end   
18'd23415: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23197;
 end   
18'd23416: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23197;
 end   
18'd23417: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23197;
 end   
18'd23418: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23197;
 end   
18'd23419: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23197;
 end   
18'd23420: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23197;
 end   
18'd23542: begin  
rid<=1;
end
18'd23543: begin  
end
18'd23544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd23545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd23546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd23547: begin  
rid<=0;
end
18'd23601: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=44;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3422;
 end   
18'd23602: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=86;
   mapp<=10;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9842;
 end   
18'd23603: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=7;
   mapp<=71;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9953;
 end   
18'd23604: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=60;
   mapp<=13;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=5727;
 end   
18'd23605: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=27;
   mapp<=15;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=13773;
 end   
18'd23606: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=85;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=9567;
 end   
18'd23607: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=18;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=14318;
 end   
18'd23608: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd23609: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd23610: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd23611: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd23612: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd23613: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=3422;
 end   
18'd23614: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=3422;
 end   
18'd23615: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=3422;
 end   
18'd23616: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=3422;
 end   
18'd23742: begin  
rid<=1;
end
18'd23743: begin  
end
18'd23744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd23745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd23746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd23747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd23748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd23749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd23750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd23751: begin  
rid<=0;
end
18'd23801: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=93;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13387;
 end   
18'd23802: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=85;
   mapp<=71;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7805;
 end   
18'd23803: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=37;
   mapp<=68;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=2997;
 end   
18'd23804: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=11;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=6122;
 end   
18'd23805: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=4;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=6123;
 end   
18'd23806: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=77;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=9104;
 end   
18'd23807: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=6;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=6696;
 end   
18'd23808: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=68;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=6052;
 end   
18'd23809: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=22;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd23810: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=13;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd23811: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd23812: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd23813: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13387;
 end   
18'd23942: begin  
rid<=1;
end
18'd23943: begin  
end
18'd23944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd23945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd23946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd23947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd23948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd23949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd23950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd23951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd23952: begin  
rid<=0;
end
18'd24001: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=93;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=17644;
 end   
18'd24002: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=84;
   mapp<=38;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=21150;
 end   
18'd24003: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=87;
   mapp<=88;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=23434;
 end   
18'd24004: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=61;
   mapp<=55;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=21651;
 end   
18'd24005: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd24006: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd24007: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd24008: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd24009: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd24010: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd24011: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd24142: begin  
rid<=1;
end
18'd24143: begin  
end
18'd24144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd24145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd24146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd24147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd24148: begin  
rid<=0;
end
18'd24201: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=82;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=82;
 end   
18'd24202: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd24342: begin  
rid<=1;
end
18'd24343: begin  
end
18'd24344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd24345: begin  
rid<=0;
end
18'd24401: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=4;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=212;
 end   
18'd24402: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=84;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4462;
 end   
18'd24403: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd24542: begin  
rid<=1;
end
18'd24543: begin  
end
18'd24544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd24545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd24546: begin  
rid<=0;
end
18'd24601: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=11;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=17687;
 end   
18'd24602: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=13;
   mapp<=64;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=17586;
 end   
18'd24603: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=68;
   mapp<=81;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=18586;
 end   
18'd24604: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=51;
   mapp<=72;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=20149;
 end   
18'd24605: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=16;
   mapp<=6;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=20725;
 end   
18'd24606: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=79;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd24607: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=68;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd24608: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd24609: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd24610: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd24611: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd24612: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd24613: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17687;
 end   
18'd24614: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17687;
 end   
18'd24615: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17687;
 end   
18'd24616: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17687;
 end   
18'd24617: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17687;
 end   
18'd24618: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17687;
 end   
18'd24742: begin  
rid<=1;
end
18'd24743: begin  
end
18'd24744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd24745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd24746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd24747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd24748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd24749: begin  
rid<=0;
end
18'd24801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=63;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6740;
 end   
18'd24802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=59;
   mapp<=79;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6144;
 end   
18'd24803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=53;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=4613;
 end   
18'd24804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=36;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=8723;
 end   
18'd24805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=95;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=8310;
 end   
18'd24806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=65;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd24807: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd24808: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd24942: begin  
rid<=1;
end
18'd24943: begin  
end
18'd24944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd24945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd24946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd24947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd24948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd24949: begin  
rid<=0;
end
18'd25001: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=8;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10521;
 end   
18'd25002: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=59;
   mapp<=80;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11432;
 end   
18'd25003: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=56;
   mapp<=76;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=11172;
 end   
18'd25004: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=2;
   mapp<=55;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=11517;
 end   
18'd25005: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=32;
   mapp<=25;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=16310;
 end   
18'd25006: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=5;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd25007: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=40;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd25008: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=75;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd25009: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd25010: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=85;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd25011: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd25012: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd25013: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10521;
 end   
18'd25014: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10521;
 end   
18'd25015: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10521;
 end   
18'd25016: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10521;
 end   
18'd25142: begin  
rid<=1;
end
18'd25143: begin  
end
18'd25144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd25145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd25146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd25147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd25148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd25149: begin  
rid<=0;
end
18'd25201: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=58;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=17477;
 end   
18'd25202: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=93;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=12782;
 end   
18'd25203: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=40;
   mapp<=2;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=11544;
 end   
18'd25204: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=46;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd25205: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=74;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd25206: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd25207: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd25208: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd25209: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd25210: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd25211: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd25212: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd25342: begin  
rid<=1;
end
18'd25343: begin  
end
18'd25344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd25345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd25346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd25347: begin  
rid<=0;
end
18'd25401: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=72;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5760;
 end   
18'd25402: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=0;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd25403: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd25404: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd25542: begin  
rid<=1;
end
18'd25543: begin  
end
18'd25544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd25545: begin  
rid<=0;
end
18'd25601: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=68;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15576;
 end   
18'd25602: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=15;
   mapp<=41;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7865;
 end   
18'd25603: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=96;
   mapp<=88;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9145;
 end   
18'd25604: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=25;
   mapp<=81;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=6021;
 end   
18'd25605: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=9;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=8749;
 end   
18'd25606: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=12;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=12180;
 end   
18'd25607: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=36;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=13630;
 end   
18'd25608: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=55;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd25609: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd25610: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=43;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd25611: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd25612: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd25613: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15576;
 end   
18'd25614: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15576;
 end   
18'd25742: begin  
rid<=1;
end
18'd25743: begin  
end
18'd25744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd25745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd25746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd25747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd25748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd25749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd25750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd25751: begin  
rid<=0;
end
18'd25801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=14;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11043;
 end   
18'd25802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=50;
   mapp<=12;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11239;
 end   
18'd25803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=90;
   mapp<=48;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=13005;
 end   
18'd25804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=35;
   mapp<=18;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=7414;
 end   
18'd25805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=59;
   mapp<=68;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=10843;
 end   
18'd25806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=69;
   mapp<=17;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=10627;
 end   
18'd25807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=95;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd25808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=3;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd25809: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=40;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd25810: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=79;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd25811: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=99;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd25812: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd25813: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11043;
 end   
18'd25814: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11043;
 end   
18'd25815: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11043;
 end   
18'd25816: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11043;
 end   
18'd25817: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11043;
 end   
18'd25942: begin  
rid<=1;
end
18'd25943: begin  
end
18'd25944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd25945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd25946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd25947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd25948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd25949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd25950: begin  
rid<=0;
end
18'd26001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=14;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=22580;
 end   
18'd26002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=18;
   mapp<=81;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=24011;
 end   
18'd26003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=44;
   mapp<=52;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=20207;
 end   
18'd26004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=63;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd26005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=29;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd26006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=52;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd26007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=64;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd26008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=69;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd26009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=70;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd26010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd26011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd26012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd26013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22580;
 end   
18'd26014: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22580;
 end   
18'd26015: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22580;
 end   
18'd26016: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22580;
 end   
18'd26017: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22580;
 end   
18'd26018: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22580;
 end   
18'd26019: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22580;
 end   
18'd26020: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22580;
 end   
18'd26142: begin  
rid<=1;
end
18'd26143: begin  
end
18'd26144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd26145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd26146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd26147: begin  
rid<=0;
end
18'd26201: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=26;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9056;
 end   
18'd26202: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=76;
   mapp<=87;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9155;
 end   
18'd26203: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=23;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5662;
 end   
18'd26204: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=40;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=10663;
 end   
18'd26205: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=79;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd26206: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd26207: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd26342: begin  
rid<=1;
end
18'd26343: begin  
end
18'd26344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd26345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd26346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd26347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd26348: begin  
rid<=0;
end
18'd26401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=62;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=21765;
 end   
18'd26402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=35;
   mapp<=71;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=27030;
 end   
18'd26403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=87;
   mapp<=45;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=28110;
 end   
18'd26404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=96;
   mapp<=21;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=30991;
 end   
18'd26405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=33;
   mapp<=70;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=30044;
 end   
18'd26406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=88;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd26407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=35;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd26408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd26409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd26410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd26411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd26412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd26413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21765;
 end   
18'd26414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21765;
 end   
18'd26415: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21765;
 end   
18'd26416: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21765;
 end   
18'd26417: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21765;
 end   
18'd26418: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21765;
 end   
18'd26542: begin  
rid<=1;
end
18'd26543: begin  
end
18'd26544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd26545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd26546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd26547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd26548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd26549: begin  
rid<=0;
end
18'd26601: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=65;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5912;
 end   
18'd26602: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=1;
   mapp<=62;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=410;
 end   
18'd26603: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=5;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=904;
 end   
18'd26604: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=7;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=4814;
 end   
18'd26605: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=67;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=10348;
 end   
18'd26606: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=69;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=8368;
 end   
18'd26607: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=34;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=7522;
 end   
18'd26608: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=71;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=9994;
 end   
18'd26609: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=57;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=11286;
 end   
18'd26610: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=98;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[9]<=11700;
 end   
18'd26611: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=45;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd26612: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd26613: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5912;
 end   
18'd26742: begin  
rid<=1;
end
18'd26743: begin  
end
18'd26744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd26745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd26746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd26747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd26748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd26749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd26750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd26751: begin  
check<=expctdoutput[7]-outcheck;
end
18'd26752: begin  
check<=expctdoutput[8]-outcheck;
end
18'd26753: begin  
check<=expctdoutput[9]-outcheck;
end
18'd26754: begin  
rid<=0;
end
18'd26801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=72;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5508;
 end   
18'd26802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=63;
   mapp<=44;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3636;
 end   
18'd26803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=28;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=3900;
 end   
18'd26804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=64;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=2506;
 end   
18'd26805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=1;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=1090;
 end   
18'd26806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=23;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=4884;
 end   
18'd26807: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=90;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd26808: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd26809: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd26942: begin  
rid<=1;
end
18'd26943: begin  
end
18'd26944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd26945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd26946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd26947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd26948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd26949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd26950: begin  
rid<=0;
end
18'd27001: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=63;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9085;
 end   
18'd27002: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=1;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=12695;
 end   
18'd27003: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=63;
   mapp<=92;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=11229;
 end   
18'd27004: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=21;
   mapp<=71;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=12029;
 end   
18'd27005: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=65;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=8682;
 end   
18'd27006: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=21;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=12647;
 end   
18'd27007: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=45;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=13896;
 end   
18'd27008: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=10;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd27009: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=95;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd27010: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=41;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd27011: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd27012: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd27013: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9085;
 end   
18'd27014: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9085;
 end   
18'd27142: begin  
rid<=1;
end
18'd27143: begin  
end
18'd27144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd27145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd27146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd27147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd27148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd27149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd27150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd27151: begin  
rid<=0;
end
18'd27201: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=54;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2754;
 end   
18'd27202: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=15;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=820;
 end   
18'd27203: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=55;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=2990;
 end   
18'd27204: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=93;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=5052;
 end   
18'd27205: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=38;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=2092;
 end   
18'd27206: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=79;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=4316;
 end   
18'd27207: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=82;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=4488;
 end   
18'd27208: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=8;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=502;
 end   
18'd27209: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd27342: begin  
rid<=1;
end
18'd27343: begin  
end
18'd27344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd27345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd27346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd27347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd27348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd27349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd27350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd27351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd27352: begin  
rid<=0;
end
18'd27401: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=4;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10110;
 end   
18'd27402: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=23;
   mapp<=38;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7762;
 end   
18'd27403: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=25;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd27404: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=78;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd27405: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=24;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd27406: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd27407: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd27408: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd27409: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd27410: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd27411: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd27542: begin  
rid<=1;
end
18'd27543: begin  
end
18'd27544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd27545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd27546: begin  
rid<=0;
end
18'd27601: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=87;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7156;
 end   
18'd27602: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=45;
   mapp<=23;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8708;
 end   
18'd27603: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=5;
   mapp<=94;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9671;
 end   
18'd27604: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=16;
   mapp<=30;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=14112;
 end   
18'd27605: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=50;
   mapp<=46;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=10809;
 end   
18'd27606: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=89;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=15295;
 end   
18'd27607: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd27608: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=63;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd27609: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=35;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd27610: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=97;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd27611: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd27612: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd27613: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7156;
 end   
18'd27614: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7156;
 end   
18'd27615: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7156;
 end   
18'd27742: begin  
rid<=1;
end
18'd27743: begin  
end
18'd27744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd27745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd27746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd27747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd27748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd27749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd27750: begin  
rid<=0;
end
18'd27801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=37;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1480;
 end   
18'd27802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=74;
   mapp<=8;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1946;
 end   
18'd27803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=20;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1076;
 end   
18'd27804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=72;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=2502;
 end   
18'd27805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=93;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd27806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd27807: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd27942: begin  
rid<=1;
end
18'd27943: begin  
end
18'd27944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd27945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd27946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd27947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd27948: begin  
rid<=0;
end
18'd28001: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=19;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3647;
 end   
18'd28002: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=41;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4008;
 end   
18'd28003: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=32;
   mapp<=6;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5978;
 end   
18'd28004: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=84;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=7325;
 end   
18'd28005: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd28006: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd28007: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd28008: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd28009: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd28142: begin  
rid<=1;
end
18'd28143: begin  
end
18'd28144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd28145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd28146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd28147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd28148: begin  
rid<=0;
end
18'd28201: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=83;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6557;
 end   
18'd28202: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=67;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5303;
 end   
18'd28203: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=36;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=2864;
 end   
18'd28204: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=25;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=2005;
 end   
18'd28205: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=18;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=1462;
 end   
18'd28206: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=37;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=2973;
 end   
18'd28207: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=28;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=2272;
 end   
18'd28208: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=19;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=1571;
 end   
18'd28209: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=77;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=6163;
 end   
18'd28210: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd28342: begin  
rid<=1;
end
18'd28343: begin  
end
18'd28344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd28345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd28346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd28347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd28348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd28349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd28350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd28351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd28352: begin  
check<=expctdoutput[8]-outcheck;
end
18'd28353: begin  
rid<=0;
end
18'd28401: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=60;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3360;
 end   
18'd28402: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=0;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=5710;
 end   
18'd28403: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd28542: begin  
rid<=1;
end
18'd28543: begin  
end
18'd28544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd28545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd28546: begin  
rid<=0;
end
18'd28601: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=36;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1152;
 end   
18'd28602: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=80;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2570;
 end   
18'd28603: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=75;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=2420;
 end   
18'd28604: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=7;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=254;
 end   
18'd28605: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=84;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=2728;
 end   
18'd28606: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd28742: begin  
rid<=1;
end
18'd28743: begin  
end
18'd28744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd28745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd28746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd28747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd28748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd28749: begin  
rid<=0;
end
18'd28801: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=51;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10484;
 end   
18'd28802: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=29;
   mapp<=76;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=12494;
 end   
18'd28803: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=90;
   mapp<=41;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=16696;
 end   
18'd28804: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=74;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=15893;
 end   
18'd28805: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=72;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=17085;
 end   
18'd28806: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=91;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=18571;
 end   
18'd28807: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd28808: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=87;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd28809: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd28810: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd28811: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd28942: begin  
rid<=1;
end
18'd28943: begin  
end
18'd28944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd28945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd28946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd28947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd28948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd28949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd28950: begin  
rid<=0;
end
18'd29001: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=39;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=20320;
 end   
18'd29002: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=68;
   mapp<=53;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=15883;
 end   
18'd29003: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=98;
   mapp<=63;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12843;
 end   
18'd29004: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=83;
   mapp<=81;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=14697;
 end   
18'd29005: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=39;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd29006: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=15;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd29007: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd29008: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd29009: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd29010: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd29011: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd29012: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd29013: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20320;
 end   
18'd29014: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20320;
 end   
18'd29015: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20320;
 end   
18'd29142: begin  
rid<=1;
end
18'd29143: begin  
end
18'd29144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd29145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd29146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd29147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd29148: begin  
rid<=0;
end
18'd29201: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=22;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=572;
 end   
18'd29202: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=38;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=998;
 end   
18'd29203: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=28;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=748;
 end   
18'd29204: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=81;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=2136;
 end   
18'd29205: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=99;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=2614;
 end   
18'd29206: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=78;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=2078;
 end   
18'd29207: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=91;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=2426;
 end   
18'd29208: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=23;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=668;
 end   
18'd29209: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd29342: begin  
rid<=1;
end
18'd29343: begin  
end
18'd29344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd29345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd29346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd29347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd29348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd29349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd29350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd29351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd29352: begin  
rid<=0;
end
18'd29401: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=41;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6829;
 end   
18'd29402: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=87;
   mapp<=49;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6472;
 end   
18'd29403: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=46;
   mapp<=2;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6622;
 end   
18'd29404: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=91;
   mapp<=7;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=5814;
 end   
18'd29405: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=37;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd29406: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=13;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd29407: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd29408: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd29409: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd29410: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd29411: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd29412: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd29413: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6829;
 end   
18'd29542: begin  
rid<=1;
end
18'd29543: begin  
end
18'd29544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd29545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd29546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd29547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd29548: begin  
rid<=0;
end
18'd29601: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=95;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=20448;
 end   
18'd29602: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=66;
   mapp<=26;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=17360;
 end   
18'd29603: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=60;
   mapp<=10;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=24469;
 end   
18'd29604: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=38;
   mapp<=77;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=23828;
 end   
18'd29605: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=88;
   mapp<=82;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=25515;
 end   
18'd29606: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=11;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd29607: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=45;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd29608: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd29609: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd29610: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd29611: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd29612: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd29613: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20448;
 end   
18'd29614: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20448;
 end   
18'd29615: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20448;
 end   
18'd29616: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20448;
 end   
18'd29617: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20448;
 end   
18'd29618: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20448;
 end   
18'd29742: begin  
rid<=1;
end
18'd29743: begin  
end
18'd29744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd29745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd29746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd29747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd29748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd29749: begin  
rid<=0;
end
18'd29801: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=23;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15896;
 end   
18'd29802: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=26;
   mapp<=89;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=18229;
 end   
18'd29803: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=3;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd29804: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=48;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd29805: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=51;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd29806: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=70;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd29807: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=36;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd29808: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=58;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd29809: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=67;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd29810: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd29811: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd29812: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd29813: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15896;
 end   
18'd29814: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15896;
 end   
18'd29815: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15896;
 end   
18'd29816: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15896;
 end   
18'd29817: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15896;
 end   
18'd29942: begin  
rid<=1;
end
18'd29943: begin  
end
18'd29944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd29945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd29946: begin  
rid<=0;
end
18'd30001: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=3;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=93;
 end   
18'd30002: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=62;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=196;
 end   
18'd30003: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=19;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=77;
 end   
18'd30004: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=75;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=255;
 end   
18'd30005: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=56;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=208;
 end   
18'd30006: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=31;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=143;
 end   
18'd30007: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=95;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=345;
 end   
18'd30008: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=44;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=202;
 end   
18'd30009: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=91;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=353;
 end   
18'd30010: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd30142: begin  
rid<=1;
end
18'd30143: begin  
end
18'd30144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd30145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd30146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd30147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd30148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd30149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd30150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd30151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd30152: begin  
check<=expctdoutput[8]-outcheck;
end
18'd30153: begin  
rid<=0;
end
18'd30201: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=19;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=950;
 end   
18'd30202: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=72;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3610;
 end   
18'd30203: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=91;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=4570;
 end   
18'd30204: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=83;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=4180;
 end   
18'd30205: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=33;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=1690;
 end   
18'd30206: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=75;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=3800;
 end   
18'd30207: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=42;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=2160;
 end   
18'd30208: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd30342: begin  
rid<=1;
end
18'd30343: begin  
end
18'd30344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd30345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd30346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd30347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd30348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd30349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd30350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd30351: begin  
rid<=0;
end
18'd30401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=50;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=23467;
 end   
18'd30402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=33;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd30403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=22;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd30404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=71;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd30405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=11;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd30406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=90;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd30407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=38;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd30408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=41;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd30409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd30410: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd30411: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd30412: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd30413: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23467;
 end   
18'd30414: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23467;
 end   
18'd30415: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23467;
 end   
18'd30416: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23467;
 end   
18'd30542: begin  
rid<=1;
end
18'd30543: begin  
end
18'd30544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd30545: begin  
rid<=0;
end
18'd30601: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=90;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=18097;
 end   
18'd30602: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=2;
   mapp<=58;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8891;
 end   
18'd30603: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=68;
   mapp<=79;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=13071;
 end   
18'd30604: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=22;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd30605: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=95;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd30606: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=35;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd30607: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=8;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd30608: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd30609: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd30610: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd30611: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd30612: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd30742: begin  
rid<=1;
end
18'd30743: begin  
end
18'd30744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd30745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd30746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd30747: begin  
rid<=0;
end
18'd30801: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=45;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4230;
 end   
18'd30802: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=99;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=4465;
 end   
18'd30803: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=88;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=3980;
 end   
18'd30804: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=78;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=3540;
 end   
18'd30805: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=42;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=1930;
 end   
18'd30806: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=57;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=2615;
 end   
18'd30807: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=41;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=1905;
 end   
18'd30808: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=47;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=2185;
 end   
18'd30809: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=69;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=3185;
 end   
18'd30810: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd30942: begin  
rid<=1;
end
18'd30943: begin  
end
18'd30944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd30945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd30946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd30947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd30948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd30949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd30950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd30951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd30952: begin  
check<=expctdoutput[8]-outcheck;
end
18'd30953: begin  
rid<=0;
end
18'd31001: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=85;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6414;
 end   
18'd31002: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=73;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd31003: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=4;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd31004: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd31005: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd31006: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd31142: begin  
rid<=1;
end
18'd31143: begin  
end
18'd31144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd31145: begin  
rid<=0;
end
18'd31201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=29;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=58;
 end   
18'd31202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=69;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=2011;
 end   
18'd31203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=54;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=1586;
 end   
18'd31204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd31342: begin  
rid<=1;
end
18'd31343: begin  
end
18'd31344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd31345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd31346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd31347: begin  
rid<=0;
end
18'd31401: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=18;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11469;
 end   
18'd31402: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=65;
   mapp<=30;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=14015;
 end   
18'd31403: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=63;
   mapp<=44;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12478;
 end   
18'd31404: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=52;
   mapp<=44;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=11515;
 end   
18'd31405: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=73;
   mapp<=49;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=9688;
 end   
18'd31406: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=70;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=10343;
 end   
18'd31407: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=31;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd31408: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=47;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd31409: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=11;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd31410: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=69;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd31411: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd31412: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd31413: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11469;
 end   
18'd31414: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11469;
 end   
18'd31415: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11469;
 end   
18'd31542: begin  
rid<=1;
end
18'd31543: begin  
end
18'd31544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd31545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd31546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd31547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd31548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd31549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd31550: begin  
rid<=0;
end
18'd31601: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=40;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14103;
 end   
18'd31602: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=11;
   mapp<=52;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11788;
 end   
18'd31603: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=92;
   mapp<=79;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=15881;
 end   
18'd31604: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=51;
   mapp<=53;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=14175;
 end   
18'd31605: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=80;
   mapp<=43;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=16031;
 end   
18'd31606: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=22;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=13428;
 end   
18'd31607: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=88;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=11711;
 end   
18'd31608: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd31609: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd31610: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd31611: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd31612: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd31613: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14103;
 end   
18'd31614: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14103;
 end   
18'd31615: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14103;
 end   
18'd31616: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14103;
 end   
18'd31742: begin  
rid<=1;
end
18'd31743: begin  
end
18'd31744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd31745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd31746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd31747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd31748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd31749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd31750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd31751: begin  
rid<=0;
end
18'd31801: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=78;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5928;
 end   
18'd31802: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=20;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1530;
 end   
18'd31803: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=15;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1160;
 end   
18'd31804: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=48;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=3678;
 end   
18'd31805: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=98;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=7488;
 end   
18'd31806: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=79;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=6054;
 end   
18'd31807: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=35;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=2720;
 end   
18'd31808: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd31942: begin  
rid<=1;
end
18'd31943: begin  
end
18'd31944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd31945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd31946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd31947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd31948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd31949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd31950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd31951: begin  
rid<=0;
end
18'd32001: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=73;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4608;
 end   
18'd32002: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=41;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2698;
 end   
18'd32003: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=62;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=5366;
 end   
18'd32004: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=20;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=4360;
 end   
18'd32005: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=70;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=6052;
 end   
18'd32006: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd32007: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd32008: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd32142: begin  
rid<=1;
end
18'd32143: begin  
end
18'd32144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd32145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd32146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd32147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd32148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd32149: begin  
rid<=0;
end
18'd32201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=67;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7952;
 end   
18'd32202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=49;
   mapp<=17;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=12027;
 end   
18'd32203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=65;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd32204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd32205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd32206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd32207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd32342: begin  
rid<=1;
end
18'd32343: begin  
end
18'd32344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd32345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd32346: begin  
rid<=0;
end
18'd32401: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=89;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5993;
 end   
18'd32402: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=52;
   mapp<=81;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8275;
 end   
18'd32403: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=30;
   mapp<=3;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=2687;
 end   
18'd32404: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=30;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=5086;
 end   
18'd32405: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd32406: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd32407: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd32408: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd32409: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd32542: begin  
rid<=1;
end
18'd32543: begin  
end
18'd32544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd32545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd32546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd32547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd32548: begin  
rid<=0;
end
18'd32601: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=40;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=32114;
 end   
18'd32602: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=33;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=34454;
 end   
18'd32603: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=37;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd32604: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=93;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd32605: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=30;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd32606: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=74;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd32607: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=93;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd32608: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=82;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd32609: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=3;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd32610: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=61;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd32611: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd32612: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd32613: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=32114;
 end   
18'd32614: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=32114;
 end   
18'd32615: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=32114;
 end   
18'd32616: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=32114;
 end   
18'd32617: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=32114;
 end   
18'd32618: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=32114;
 end   
18'd32619: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=32114;
 end   
18'd32620: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=32114;
 end   
18'd32621: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=32114;
 end   
18'd32742: begin  
rid<=1;
end
18'd32743: begin  
end
18'd32744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd32745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd32746: begin  
rid<=0;
end
18'd32801: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=66;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=18493;
 end   
18'd32802: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=83;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=21563;
 end   
18'd32803: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=61;
   mapp<=51;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=13846;
 end   
18'd32804: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=59;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd32805: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=45;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd32806: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=86;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd32807: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd32808: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd32809: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd32810: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd32811: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd32812: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd32813: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18493;
 end   
18'd32814: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18493;
 end   
18'd32942: begin  
rid<=1;
end
18'd32943: begin  
end
18'd32944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd32945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd32946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd32947: begin  
rid<=0;
end
18'd33001: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=83;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4642;
 end   
18'd33002: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=50;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9844;
 end   
18'd33003: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=58;
   mapp<=9;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9450;
 end   
18'd33004: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=21;
   mapp<=97;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=12219;
 end   
18'd33005: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=75;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=11025;
 end   
18'd33006: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=81;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd33007: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=87;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd33008: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=71;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd33009: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd33010: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd33011: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd33012: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd33142: begin  
rid<=1;
end
18'd33143: begin  
end
18'd33144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd33145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd33146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd33147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd33148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd33149: begin  
rid<=0;
end
18'd33201: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=28;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7409;
 end   
18'd33202: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=59;
   mapp<=79;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11064;
 end   
18'd33203: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=22;
   mapp<=38;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8802;
 end   
18'd33204: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=98;
   mapp<=0;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=5206;
 end   
18'd33205: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=60;
   mapp<=30;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=7765;
 end   
18'd33206: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd33207: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd33208: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd33209: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd33210: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd33211: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd33212: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd33213: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7409;
 end   
18'd33214: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7409;
 end   
18'd33342: begin  
rid<=1;
end
18'd33343: begin  
end
18'd33344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd33345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd33346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd33347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd33348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd33349: begin  
rid<=0;
end
18'd33401: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=46;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=23133;
 end   
18'd33402: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=38;
   mapp<=14;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=19999;
 end   
18'd33403: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=70;
   mapp<=67;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=22392;
 end   
18'd33404: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=38;
   mapp<=93;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=19914;
 end   
18'd33405: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=76;
   mapp<=96;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=23640;
 end   
18'd33406: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=55;
   mapp<=61;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=23610;
 end   
18'd33407: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=17;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd33408: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=71;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd33409: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=60;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd33410: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=52;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd33411: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=58;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd33412: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd33413: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23133;
 end   
18'd33414: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23133;
 end   
18'd33415: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23133;
 end   
18'd33416: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23133;
 end   
18'd33417: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23133;
 end   
18'd33542: begin  
rid<=1;
end
18'd33543: begin  
end
18'd33544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd33545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd33546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd33547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd33548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd33549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd33550: begin  
rid<=0;
end
18'd33601: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=26;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1690;
 end   
18'd33602: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=1;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=75;
 end   
18'd33603: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=34;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=2230;
 end   
18'd33604: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=59;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=3865;
 end   
18'd33605: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd33742: begin  
rid<=1;
end
18'd33743: begin  
end
18'd33744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd33745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd33746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd33747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd33748: begin  
rid<=0;
end
18'd33801: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=27;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10987;
 end   
18'd33802: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=98;
   mapp<=92;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11608;
 end   
18'd33803: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=93;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=5765;
 end   
18'd33804: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=33;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=4547;
 end   
18'd33805: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=37;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=1333;
 end   
18'd33806: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=3;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=8951;
 end   
18'd33807: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=90;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=3568;
 end   
18'd33808: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=11;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=9579;
 end   
18'd33809: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=94;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=9282;
 end   
18'd33810: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd33811: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd33812: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd33942: begin  
rid<=1;
end
18'd33943: begin  
end
18'd33944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd33945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd33946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd33947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd33948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd33949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd33950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd33951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd33952: begin  
check<=expctdoutput[8]-outcheck;
end
18'd33953: begin  
rid<=0;
end
18'd34001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=43;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7500;
 end   
18'd34002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=31;
   mapp<=47;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5224;
 end   
18'd34003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=54;
   mapp<=49;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6814;
 end   
18'd34004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=31;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=7552;
 end   
18'd34005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=69;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=10624;
 end   
18'd34006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=75;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=8959;
 end   
18'd34007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=98;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=7737;
 end   
18'd34008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=49;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=8639;
 end   
18'd34009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=36;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=5939;
 end   
18'd34010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd34011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd34012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd34013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7500;
 end   
18'd34014: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7500;
 end   
18'd34142: begin  
rid<=1;
end
18'd34143: begin  
end
18'd34144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd34145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd34146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd34147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd34148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd34149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd34150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd34151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd34152: begin  
check<=expctdoutput[8]-outcheck;
end
18'd34153: begin  
rid<=0;
end
18'd34201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=4;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4762;
 end   
18'd34202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=66;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1334;
 end   
18'd34203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=16;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=6222;
 end   
18'd34204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd34205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd34206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd34342: begin  
rid<=1;
end
18'd34343: begin  
end
18'd34344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd34345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd34346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd34347: begin  
rid<=0;
end
18'd34401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=43;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15391;
 end   
18'd34402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=4;
   mapp<=84;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=14175;
 end   
18'd34403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=99;
   mapp<=92;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=14102;
 end   
18'd34404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=74;
   mapp<=67;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=12154;
 end   
18'd34405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=48;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=6164;
 end   
18'd34406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=69;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=5262;
 end   
18'd34407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=30;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=9440;
 end   
18'd34408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=11;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=11507;
 end   
18'd34409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd34410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd34411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd34412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd34413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15391;
 end   
18'd34414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15391;
 end   
18'd34415: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15391;
 end   
18'd34542: begin  
rid<=1;
end
18'd34543: begin  
end
18'd34544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd34545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd34546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd34547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd34548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd34549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd34550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd34551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd34552: begin  
rid<=0;
end
18'd34601: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=58;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3364;
 end   
18'd34602: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=0;
   mapp<=89;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=5172;
 end   
18'd34603: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd34742: begin  
rid<=1;
end
18'd34743: begin  
end
18'd34744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd34745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd34746: begin  
rid<=0;
end
18'd34801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=18;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3406;
 end   
18'd34802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=64;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6018;
 end   
18'd34803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=75;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=4585;
 end   
18'd34804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=26;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd34805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd34806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd34942: begin  
rid<=1;
end
18'd34943: begin  
end
18'd34944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd34945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd34946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd34947: begin  
rid<=0;
end
18'd35001: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=87;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=30663;
 end   
18'd35002: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=83;
   mapp<=12;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=30170;
 end   
18'd35003: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=85;
   mapp<=40;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=36571;
 end   
18'd35004: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=90;
   mapp<=70;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=33374;
 end   
18'd35005: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=50;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd35006: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=86;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd35007: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=55;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd35008: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd35009: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd35010: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd35011: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd35012: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd35013: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=30663;
 end   
18'd35014: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=30663;
 end   
18'd35015: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=30663;
 end   
18'd35016: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=30663;
 end   
18'd35017: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=30663;
 end   
18'd35142: begin  
rid<=1;
end
18'd35143: begin  
end
18'd35144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd35145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd35146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd35147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd35148: begin  
rid<=0;
end
18'd35201: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=28;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3598;
 end   
18'd35202: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=46;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5018;
 end   
18'd35203: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=62;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=2860;
 end   
18'd35204: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=24;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=3692;
 end   
18'd35205: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=65;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=5172;
 end   
18'd35206: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=72;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=3538;
 end   
18'd35207: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=32;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=4866;
 end   
18'd35208: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd35209: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd35210: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd35342: begin  
rid<=1;
end
18'd35343: begin  
end
18'd35344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd35345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd35346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd35347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd35348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd35349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd35350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd35351: begin  
rid<=0;
end
18'd35401: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=25;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2075;
 end   
18'd35402: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=65;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5405;
 end   
18'd35403: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=60;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5000;
 end   
18'd35404: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=45;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=3765;
 end   
18'd35405: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=78;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=6514;
 end   
18'd35406: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=21;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=1793;
 end   
18'd35407: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=55;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=4625;
 end   
18'd35408: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=20;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=1730;
 end   
18'd35409: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=27;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=2321;
 end   
18'd35410: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=73;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[9]<=6149;
 end   
18'd35411: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=34;
   mapp<=0;
   pp<=100;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[10]<=2922;
 end   
18'd35412: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd35542: begin  
rid<=1;
end
18'd35543: begin  
end
18'd35544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd35545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd35546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd35547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd35548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd35549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd35550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd35551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd35552: begin  
check<=expctdoutput[8]-outcheck;
end
18'd35553: begin  
check<=expctdoutput[9]-outcheck;
end
18'd35554: begin  
check<=expctdoutput[10]-outcheck;
end
18'd35555: begin  
rid<=0;
end
18'd35601: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=74;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9207;
 end   
18'd35602: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=90;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd35603: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=56;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd35604: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=71;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd35605: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=80;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd35606: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd35607: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd35608: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd35609: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd35610: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd35742: begin  
rid<=1;
end
18'd35743: begin  
end
18'd35744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd35745: begin  
rid<=0;
end
18'd35801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=18;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3301;
 end   
18'd35802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=73;
   mapp<=25;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6296;
 end   
18'd35803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=12;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1929;
 end   
18'd35804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd35805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd35806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd35942: begin  
rid<=1;
end
18'd35943: begin  
end
18'd35944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd35945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd35946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd35947: begin  
rid<=0;
end
18'd36001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=46;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8173;
 end   
18'd36002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=3;
   mapp<=17;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6350;
 end   
18'd36003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=31;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd36004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=15;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd36005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=39;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd36006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=58;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd36007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd36008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd36009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd36010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd36011: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd36142: begin  
rid<=1;
end
18'd36143: begin  
end
18'd36144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd36145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd36146: begin  
rid<=0;
end
18'd36201: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=73;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=27122;
 end   
18'd36202: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=80;
   mapp<=99;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=24028;
 end   
18'd36203: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=38;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd36204: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=97;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd36205: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=42;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd36206: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=8;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd36207: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd36208: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd36209: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd36210: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd36211: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd36212: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd36213: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=27122;
 end   
18'd36342: begin  
rid<=1;
end
18'd36343: begin  
end
18'd36344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd36345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd36346: begin  
rid<=0;
end
18'd36401: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=38;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1664;
 end   
18'd36402: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=21;
   mapp<=34;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1323;
 end   
18'd36403: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=1;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=1696;
 end   
18'd36404: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=78;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=4716;
 end   
18'd36405: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=82;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=4605;
 end   
18'd36406: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=69;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=3428;
 end   
18'd36407: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=36;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=3066;
 end   
18'd36408: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=78;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=3853;
 end   
18'd36409: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd36410: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd36411: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd36542: begin  
rid<=1;
end
18'd36543: begin  
end
18'd36544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd36545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd36546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd36547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd36548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd36549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd36550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd36551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd36552: begin  
rid<=0;
end
18'd36601: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=16;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11708;
 end   
18'd36602: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=37;
   mapp<=75;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7789;
 end   
18'd36603: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=7;
   mapp<=24;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=14282;
 end   
18'd36604: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=93;
   mapp<=81;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=7687;
 end   
18'd36605: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=84;
   mapp<=0;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=6949;
 end   
18'd36606: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=61;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=15778;
 end   
18'd36607: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=62;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=17353;
 end   
18'd36608: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd36609: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd36610: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd36611: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd36612: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd36613: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11708;
 end   
18'd36614: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11708;
 end   
18'd36615: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11708;
 end   
18'd36616: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11708;
 end   
18'd36742: begin  
rid<=1;
end
18'd36743: begin  
end
18'd36744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd36745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd36746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd36747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd36748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd36749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd36750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd36751: begin  
rid<=0;
end
18'd36801: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=91;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16679;
 end   
18'd36802: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=64;
   mapp<=58;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=12711;
 end   
18'd36803: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=23;
   mapp<=43;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12214;
 end   
18'd36804: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=15;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd36805: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=72;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd36806: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=29;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd36807: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=41;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd36808: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=15;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd36809: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=15;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd36810: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=36;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd36811: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd36812: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd36813: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16679;
 end   
18'd36814: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16679;
 end   
18'd36815: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16679;
 end   
18'd36816: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16679;
 end   
18'd36817: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16679;
 end   
18'd36818: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16679;
 end   
18'd36942: begin  
rid<=1;
end
18'd36943: begin  
end
18'd36944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd36945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd36946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd36947: begin  
rid<=0;
end
18'd37001: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=24;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16538;
 end   
18'd37002: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=74;
   mapp<=52;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=21748;
 end   
18'd37003: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=33;
   mapp<=93;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=19697;
 end   
18'd37004: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=85;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd37005: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=38;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd37006: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=70;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd37007: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=62;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd37008: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd37009: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd37010: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd37011: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd37012: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd37013: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16538;
 end   
18'd37014: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16538;
 end   
18'd37015: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16538;
 end   
18'd37016: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16538;
 end   
18'd37142: begin  
rid<=1;
end
18'd37143: begin  
end
18'd37144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd37145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd37146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd37147: begin  
rid<=0;
end
18'd37201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4011;
 end   
18'd37202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=24;
   mapp<=78;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8467;
 end   
18'd37203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=93;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd37204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd37205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd37206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd37207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd37342: begin  
rid<=1;
end
18'd37343: begin  
end
18'd37344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd37345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd37346: begin  
rid<=0;
end
18'd37401: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=90;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=17658;
 end   
18'd37402: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=34;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=18225;
 end   
18'd37403: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=91;
   mapp<=7;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=18283;
 end   
18'd37404: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=21;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd37405: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=85;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd37406: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=34;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd37407: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=90;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd37408: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=42;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd37409: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd37410: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd37411: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd37412: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd37413: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17658;
 end   
18'd37414: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17658;
 end   
18'd37542: begin  
rid<=1;
end
18'd37543: begin  
end
18'd37544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd37545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd37546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd37547: begin  
rid<=0;
end
18'd37601: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=97;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4638;
 end   
18'd37602: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=76;
   mapp<=21;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4168;
 end   
18'd37603: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=54;
   mapp<=24;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=2633;
 end   
18'd37604: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=69;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=2088;
 end   
18'd37605: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=8;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=2983;
 end   
18'd37606: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=27;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=4121;
 end   
18'd37607: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=93;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=4746;
 end   
18'd37608: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=68;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=2728;
 end   
18'd37609: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=66;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd37610: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=2;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd37611: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd37612: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd37613: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=4638;
 end   
18'd37742: begin  
rid<=1;
end
18'd37743: begin  
end
18'd37744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd37745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd37746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd37747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd37748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd37749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd37750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd37751: begin  
check<=expctdoutput[7]-outcheck;
end
18'd37752: begin  
rid<=0;
end
18'd37801: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=78;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16846;
 end   
18'd37802: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=14;
   mapp<=18;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=15807;
 end   
18'd37803: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=87;
   mapp<=90;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=15025;
 end   
18'd37804: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=39;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd37805: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=74;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd37806: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=20;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd37807: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd37808: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd37809: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd37810: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd37811: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd37812: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd37813: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16846;
 end   
18'd37814: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16846;
 end   
18'd37942: begin  
rid<=1;
end
18'd37943: begin  
end
18'd37944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd37945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd37946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd37947: begin  
rid<=0;
end
18'd38001: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=2;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1429;
 end   
18'd38002: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=21;
   mapp<=41;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2318;
 end   
18'd38003: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=4;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd38004: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd38005: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd38006: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd38007: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd38142: begin  
rid<=1;
end
18'd38143: begin  
end
18'd38144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd38145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd38146: begin  
rid<=0;
end
18'd38201: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=60;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15392;
 end   
18'd38202: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=61;
   mapp<=33;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=12173;
 end   
18'd38203: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=20;
   mapp<=8;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=16286;
 end   
18'd38204: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=43;
   mapp<=61;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=17879;
 end   
18'd38205: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=78;
   mapp<=33;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=17931;
 end   
18'd38206: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=87;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd38207: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd38208: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd38209: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd38210: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd38211: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd38212: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd38213: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15392;
 end   
18'd38214: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15392;
 end   
18'd38215: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15392;
 end   
18'd38216: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15392;
 end   
18'd38342: begin  
rid<=1;
end
18'd38343: begin  
end
18'd38344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd38345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd38346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd38347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd38348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd38349: begin  
rid<=0;
end
18'd38401: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=61;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9428;
 end   
18'd38402: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=12;
   mapp<=34;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5217;
 end   
18'd38403: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=11;
   mapp<=15;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5920;
 end   
18'd38404: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=59;
   mapp<=56;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=11623;
 end   
18'd38405: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=51;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd38406: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd38407: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd38408: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd38409: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd38410: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd38411: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd38542: begin  
rid<=1;
end
18'd38543: begin  
end
18'd38544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd38545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd38546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd38547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd38548: begin  
rid<=0;
end
18'd38601: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=60;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=30097;
 end   
18'd38602: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=93;
   mapp<=84;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=23642;
 end   
18'd38603: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=72;
   mapp<=51;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=18424;
 end   
18'd38604: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=2;
   mapp<=1;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=24530;
 end   
18'd38605: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=76;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd38606: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=43;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd38607: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=73;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd38608: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=66;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd38609: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd38610: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd38611: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd38612: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd38613: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=30097;
 end   
18'd38614: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=30097;
 end   
18'd38615: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=30097;
 end   
18'd38616: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=30097;
 end   
18'd38617: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=30097;
 end   
18'd38618: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=30097;
 end   
18'd38619: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=30097;
 end   
18'd38742: begin  
rid<=1;
end
18'd38743: begin  
end
18'd38744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd38745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd38746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd38747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd38748: begin  
rid<=0;
end
18'd38801: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=53;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11546;
 end   
18'd38802: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=92;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=23245;
 end   
18'd38803: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=70;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd38804: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=19;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd38805: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=72;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd38806: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=7;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd38807: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=94;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd38808: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=5;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd38809: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd38810: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd38811: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd38812: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd38813: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11546;
 end   
18'd38814: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11546;
 end   
18'd38815: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11546;
 end   
18'd38816: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11546;
 end   
18'd38817: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11546;
 end   
18'd38942: begin  
rid<=1;
end
18'd38943: begin  
end
18'd38944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd38945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd38946: begin  
rid<=0;
end
18'd39001: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=71;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4402;
 end   
18'd39002: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=9;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=649;
 end   
18'd39003: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=7;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=517;
 end   
18'd39004: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=38;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=2728;
 end   
18'd39005: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=60;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=4300;
 end   
18'd39006: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=71;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=5091;
 end   
18'd39007: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd39142: begin  
rid<=1;
end
18'd39143: begin  
end
18'd39144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd39145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd39146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd39147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd39148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd39149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd39150: begin  
rid<=0;
end
18'd39201: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=70;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16447;
 end   
18'd39202: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=39;
   mapp<=23;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=20658;
 end   
18'd39203: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=66;
   mapp<=29;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=18359;
 end   
18'd39204: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=22;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd39205: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=83;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd39206: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=60;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd39207: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd39208: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd39209: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd39210: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd39211: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd39212: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd39213: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16447;
 end   
18'd39214: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16447;
 end   
18'd39342: begin  
rid<=1;
end
18'd39343: begin  
end
18'd39344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd39345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd39346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd39347: begin  
rid<=0;
end
18'd39401: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=88;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=28785;
 end   
18'd39402: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=52;
   mapp<=59;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=25002;
 end   
18'd39403: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=54;
   mapp<=86;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=26656;
 end   
18'd39404: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=66;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd39405: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=33;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd39406: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=60;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd39407: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=19;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd39408: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=31;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd39409: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=38;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd39410: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=67;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd39411: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=76;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd39412: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd39413: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28785;
 end   
18'd39414: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28785;
 end   
18'd39415: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28785;
 end   
18'd39416: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28785;
 end   
18'd39417: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28785;
 end   
18'd39418: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28785;
 end   
18'd39419: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28785;
 end   
18'd39420: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28785;
 end   
18'd39542: begin  
rid<=1;
end
18'd39543: begin  
end
18'd39544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd39545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd39546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd39547: begin  
rid<=0;
end
18'd39601: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=53;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1060;
 end   
18'd39602: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=7;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=150;
 end   
18'd39603: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=69;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1400;
 end   
18'd39604: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=16;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=350;
 end   
18'd39605: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=22;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=480;
 end   
18'd39606: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd39742: begin  
rid<=1;
end
18'd39743: begin  
end
18'd39744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd39745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd39746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd39747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd39748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd39749: begin  
rid<=0;
end
18'd39801: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=17;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1071;
 end   
18'd39802: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=60;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=1030;
 end   
18'd39803: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=47;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=819;
 end   
18'd39804: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=93;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=1611;
 end   
18'd39805: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=30;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=550;
 end   
18'd39806: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=17;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=339;
 end   
18'd39807: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=43;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=791;
 end   
18'd39808: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=76;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=1362;
 end   
18'd39809: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=14;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=318;
 end   
18'd39810: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=26;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[9]<=532;
 end   
18'd39811: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd39942: begin  
rid<=1;
end
18'd39943: begin  
end
18'd39944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd39945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd39946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd39947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd39948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd39949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd39950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd39951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd39952: begin  
check<=expctdoutput[8]-outcheck;
end
18'd39953: begin  
check<=expctdoutput[9]-outcheck;
end
18'd39954: begin  
rid<=0;
end
18'd40001: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=66;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=21388;
 end   
18'd40002: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=93;
   mapp<=92;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=17301;
 end   
18'd40003: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=64;
   mapp<=64;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12112;
 end   
18'd40004: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=75;
   mapp<=54;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=6123;
 end   
18'd40005: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd40006: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd40007: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd40008: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd40009: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd40010: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd40011: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd40142: begin  
rid<=1;
end
18'd40143: begin  
end
18'd40144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd40145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd40146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd40147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd40148: begin  
rid<=0;
end
18'd40201: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=72;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5688;
 end   
18'd40202: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=43;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=3106;
 end   
18'd40203: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=77;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=5564;
 end   
18'd40204: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=89;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=6438;
 end   
18'd40205: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=61;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=4432;
 end   
18'd40206: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=85;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=6170;
 end   
18'd40207: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd40342: begin  
rid<=1;
end
18'd40343: begin  
end
18'd40344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd40345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd40346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd40347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd40348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd40349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd40350: begin  
rid<=0;
end
18'd40401: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=57;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15283;
 end   
18'd40402: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=30;
   mapp<=63;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11293;
 end   
18'd40403: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=23;
   mapp<=4;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=11771;
 end   
18'd40404: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=64;
   mapp<=46;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=17754;
 end   
18'd40405: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=74;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd40406: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=46;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd40407: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd40408: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=81;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd40409: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=18;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd40410: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd40411: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd40412: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd40413: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15283;
 end   
18'd40414: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15283;
 end   
18'd40415: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15283;
 end   
18'd40542: begin  
rid<=1;
end
18'd40543: begin  
end
18'd40544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd40545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd40546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd40547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd40548: begin  
rid<=0;
end
18'd40601: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=61;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8463;
 end   
18'd40602: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=91;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4055;
 end   
18'd40603: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd40604: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd40605: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd40742: begin  
rid<=1;
end
18'd40743: begin  
end
18'd40744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd40745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd40746: begin  
rid<=0;
end
18'd40801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=91;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8918;
 end   
18'd40802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=0;
   mapp<=69;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5461;
 end   
18'd40803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=79;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8935;
 end   
18'd40804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=17;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=2869;
 end   
18'd40805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=17;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=2672;
 end   
18'd40806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=14;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=7977;
 end   
18'd40807: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=95;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd40808: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd40809: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd40942: begin  
rid<=1;
end
18'd40943: begin  
end
18'd40944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd40945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd40946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd40947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd40948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd40949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd40950: begin  
rid<=0;
end
18'd41001: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=28;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1876;
 end   
18'd41002: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=53;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3561;
 end   
18'd41003: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=9;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=623;
 end   
18'd41004: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=73;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=4921;
 end   
18'd41005: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=81;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=5467;
 end   
18'd41006: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=3;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=251;
 end   
18'd41007: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=69;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=4683;
 end   
18'd41008: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=16;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=1142;
 end   
18'd41009: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd41142: begin  
rid<=1;
end
18'd41143: begin  
end
18'd41144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd41145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd41146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd41147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd41148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd41149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd41150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd41151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd41152: begin  
rid<=0;
end
18'd41201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=57;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5007;
 end   
18'd41202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=81;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2554;
 end   
18'd41203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd41204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd41205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd41342: begin  
rid<=1;
end
18'd41343: begin  
end
18'd41344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd41345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd41346: begin  
rid<=0;
end
18'd41401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=77;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13541;
 end   
18'd41402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=45;
   mapp<=87;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11246;
 end   
18'd41403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=64;
   mapp<=71;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12591;
 end   
18'd41404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=38;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=12052;
 end   
18'd41405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=71;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd41406: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=47;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd41407: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd41408: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd41409: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd41542: begin  
rid<=1;
end
18'd41543: begin  
end
18'd41544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd41545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd41546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd41547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd41548: begin  
rid<=0;
end
18'd41601: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=5;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3076;
 end   
18'd41602: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=53;
   mapp<=57;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4640;
 end   
18'd41603: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=71;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5361;
 end   
18'd41604: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=80;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=3190;
 end   
18'd41605: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=40;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=2190;
 end   
18'd41606: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=30;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd41607: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd41608: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd41742: begin  
rid<=1;
end
18'd41743: begin  
end
18'd41744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd41745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd41746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd41747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd41748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd41749: begin  
rid<=0;
end
18'd41801: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=86;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16770;
 end   
18'd41802: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=4;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10261;
 end   
18'd41803: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=89;
   mapp<=98;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=14729;
 end   
18'd41804: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=31;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=14832;
 end   
18'd41805: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=44;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=11756;
 end   
18'd41806: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=88;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=10504;
 end   
18'd41807: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=10;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=4208;
 end   
18'd41808: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=18;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=8935;
 end   
18'd41809: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=19;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=8979;
 end   
18'd41810: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=59;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd41811: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=27;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd41812: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd41813: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16770;
 end   
18'd41814: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16770;
 end   
18'd41942: begin  
rid<=1;
end
18'd41943: begin  
end
18'd41944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd41945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd41946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd41947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd41948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd41949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd41950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd41951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd41952: begin  
check<=expctdoutput[8]-outcheck;
end
18'd41953: begin  
rid<=0;
end
18'd42001: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=0;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1536;
 end   
18'd42002: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=96;
   mapp<=16;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8442;
 end   
18'd42003: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=53;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5135;
 end   
18'd42004: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=58;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd42005: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd42006: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd42142: begin  
rid<=1;
end
18'd42143: begin  
end
18'd42144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd42145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd42146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd42147: begin  
rid<=0;
end
18'd42201: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=46;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=18979;
 end   
18'd42202: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=29;
   mapp<=49;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=20787;
 end   
18'd42203: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=71;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd42204: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=28;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd42205: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=59;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd42206: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=41;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd42207: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=21;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd42208: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=88;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd42209: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=66;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd42210: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd42211: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd42212: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd42213: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18979;
 end   
18'd42214: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18979;
 end   
18'd42215: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18979;
 end   
18'd42216: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18979;
 end   
18'd42217: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18979;
 end   
18'd42342: begin  
rid<=1;
end
18'd42343: begin  
end
18'd42344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd42345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd42346: begin  
rid<=0;
end
18'd42401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=87;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=35635;
 end   
18'd42402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=38;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd42403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=69;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd42404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=83;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd42405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=40;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd42406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=95;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd42407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=66;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd42408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=33;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd42409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=9;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd42410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=57;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd42411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=17;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd42412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd42413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=35635;
 end   
18'd42414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=35635;
 end   
18'd42415: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=35635;
 end   
18'd42416: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=35635;
 end   
18'd42417: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=35635;
 end   
18'd42418: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=35635;
 end   
18'd42419: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=35635;
 end   
18'd42420: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=35635;
 end   
18'd42421: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=35635;
 end   
18'd42422: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=35635;
 end   
18'd42542: begin  
rid<=1;
end
18'd42543: begin  
end
18'd42544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd42545: begin  
rid<=0;
end
18'd42601: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=74;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=37417;
 end   
18'd42602: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=12;
   mapp<=58;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=32010;
 end   
18'd42603: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=97;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd42604: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=51;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd42605: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=95;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd42606: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=17;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd42607: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=92;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd42608: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=92;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd42609: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=37;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd42610: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=30;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd42611: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=13;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd42612: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd42613: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=37417;
 end   
18'd42614: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=37417;
 end   
18'd42615: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=37417;
 end   
18'd42616: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=37417;
 end   
18'd42617: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=37417;
 end   
18'd42618: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=37417;
 end   
18'd42619: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=37417;
 end   
18'd42620: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=37417;
 end   
18'd42621: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=37417;
 end   
18'd42742: begin  
rid<=1;
end
18'd42743: begin  
end
18'd42744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd42745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd42746: begin  
rid<=0;
end
18'd42801: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=20;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=19300;
 end   
18'd42802: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=93;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd42803: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=92;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd42804: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=62;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd42805: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=14;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd42806: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=27;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd42807: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=7;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd42808: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=94;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd42809: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd42810: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd42811: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd42812: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd42813: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19300;
 end   
18'd42814: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19300;
 end   
18'd42815: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19300;
 end   
18'd42816: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19300;
 end   
18'd42942: begin  
rid<=1;
end
18'd42943: begin  
end
18'd42944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd42945: begin  
rid<=0;
end
18'd43001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=95;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12355;
 end   
18'd43002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=62;
   mapp<=13;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6743;
 end   
18'd43003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=81;
   mapp<=93;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5622;
 end   
18'd43004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=46;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd43005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=9;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd43006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=48;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd43007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=68;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd43008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd43009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd43010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd43011: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd43012: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd43142: begin  
rid<=1;
end
18'd43143: begin  
end
18'd43144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd43145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd43146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd43147: begin  
rid<=0;
end
18'd43201: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=62;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8533;
 end   
18'd43202: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=27;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7622;
 end   
18'd43203: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=77;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd43204: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=17;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd43205: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=40;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd43206: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=42;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd43207: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd43208: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd43209: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd43210: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd43211: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd43342: begin  
rid<=1;
end
18'd43343: begin  
end
18'd43344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd43345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd43346: begin  
rid<=0;
end
18'd43401: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=22;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=18983;
 end   
18'd43402: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=27;
   mapp<=76;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=17818;
 end   
18'd43403: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=29;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd43404: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=11;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd43405: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=11;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd43406: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=54;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd43407: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=80;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd43408: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=53;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd43409: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=93;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd43410: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=21;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd43411: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd43412: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd43413: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18983;
 end   
18'd43414: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18983;
 end   
18'd43415: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18983;
 end   
18'd43416: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18983;
 end   
18'd43417: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18983;
 end   
18'd43418: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18983;
 end   
18'd43419: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18983;
 end   
18'd43542: begin  
rid<=1;
end
18'd43543: begin  
end
18'd43544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd43545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd43546: begin  
rid<=0;
end
18'd43601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=31;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=17431;
 end   
18'd43602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=40;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=17837;
 end   
18'd43603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=34;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd43604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=40;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd43605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=86;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd43606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=34;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd43607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=48;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd43608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=39;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd43609: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd43610: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd43611: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd43612: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd43613: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17431;
 end   
18'd43614: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17431;
 end   
18'd43615: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17431;
 end   
18'd43742: begin  
rid<=1;
end
18'd43743: begin  
end
18'd43744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd43745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd43746: begin  
rid<=0;
end
18'd43801: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=62;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=744;
 end   
18'd43802: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=52;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=634;
 end   
18'd43803: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=31;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=392;
 end   
18'd43804: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=87;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=1074;
 end   
18'd43805: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd43942: begin  
rid<=1;
end
18'd43943: begin  
end
18'd43944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd43945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd43946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd43947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd43948: begin  
rid<=0;
end
18'd44001: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=56;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2688;
 end   
18'd44002: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=70;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3370;
 end   
18'd44003: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=50;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=2420;
 end   
18'd44004: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=82;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=3966;
 end   
18'd44005: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=1;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=88;
 end   
18'd44006: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=93;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=4514;
 end   
18'd44007: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=99;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=4812;
 end   
18'd44008: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=32;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=1606;
 end   
18'd44009: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=44;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=2192;
 end   
18'd44010: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd44142: begin  
rid<=1;
end
18'd44143: begin  
end
18'd44144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd44145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd44146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd44147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd44148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd44149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd44150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd44151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd44152: begin  
check<=expctdoutput[8]-outcheck;
end
18'd44153: begin  
rid<=0;
end
18'd44201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=66;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2190;
 end   
18'd44202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=38;
   mapp<=50;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=810;
 end   
18'd44203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=1;
   mapp<=26;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=2292;
 end   
18'd44204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=23;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=3338;
 end   
18'd44205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=43;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=4342;
 end   
18'd44206: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=41;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=6684;
 end   
18'd44207: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=80;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=5598;
 end   
18'd44208: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=95;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=2884;
 end   
18'd44209: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=18;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd44210: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=59;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd44211: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd44212: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd44213: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=2190;
 end   
18'd44342: begin  
rid<=1;
end
18'd44343: begin  
end
18'd44344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd44345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd44346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd44347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd44348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd44349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd44350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd44351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd44352: begin  
rid<=0;
end
18'd44401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=15;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=435;
 end   
18'd44402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=88;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=1330;
 end   
18'd44403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=54;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=830;
 end   
18'd44404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=13;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=225;
 end   
18'd44405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=79;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=1225;
 end   
18'd44406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=69;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=1085;
 end   
18'd44407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=66;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=1050;
 end   
18'd44408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=79;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=1255;
 end   
18'd44409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=77;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=1235;
 end   
18'd44410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=37;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[9]<=645;
 end   
18'd44411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=2;
   pp<=100;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[10]<=130;
 end   
18'd44412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd44542: begin  
rid<=1;
end
18'd44543: begin  
end
18'd44544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd44545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd44546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd44547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd44548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd44549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd44550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd44551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd44552: begin  
check<=expctdoutput[8]-outcheck;
end
18'd44553: begin  
check<=expctdoutput[9]-outcheck;
end
18'd44554: begin  
check<=expctdoutput[10]-outcheck;
end
18'd44555: begin  
rid<=0;
end
18'd44601: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=97;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=18774;
 end   
18'd44602: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=8;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=16967;
 end   
18'd44603: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=8;
   mapp<=23;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=10786;
 end   
18'd44604: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=11;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd44605: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=93;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd44606: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=65;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd44607: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=81;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd44608: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=2;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd44609: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd44610: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd44611: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd44612: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd44613: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18774;
 end   
18'd44614: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18774;
 end   
18'd44742: begin  
rid<=1;
end
18'd44743: begin  
end
18'd44744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd44745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd44746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd44747: begin  
rid<=0;
end
18'd44801: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=40;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2405;
 end   
18'd44802: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=33;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2355;
 end   
18'd44803: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=65;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=3379;
 end   
18'd44804: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=23;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=3227;
 end   
18'd44805: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=69;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=3295;
 end   
18'd44806: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=15;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=2399;
 end   
18'd44807: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=53;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=2345;
 end   
18'd44808: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=5;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=3042;
 end   
18'd44809: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=84;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=6014;
 end   
18'd44810: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=78;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[9]<=4695;
 end   
18'd44811: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd44812: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd44813: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=2405;
 end   
18'd44942: begin  
rid<=1;
end
18'd44943: begin  
end
18'd44944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd44945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd44946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd44947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd44948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd44949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd44950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd44951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd44952: begin  
check<=expctdoutput[8]-outcheck;
end
18'd44953: begin  
check<=expctdoutput[9]-outcheck;
end
18'd44954: begin  
rid<=0;
end
18'd45001: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=85;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12965;
 end   
18'd45002: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=48;
   mapp<=94;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11944;
 end   
18'd45003: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=81;
   mapp<=33;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=10384;
 end   
18'd45004: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=32;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=7800;
 end   
18'd45005: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=56;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd45006: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=10;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd45007: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd45008: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd45009: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd45142: begin  
rid<=1;
end
18'd45143: begin  
end
18'd45144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd45145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd45146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd45147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd45148: begin  
rid<=0;
end
18'd45201: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=27;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8177;
 end   
18'd45202: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=37;
   mapp<=6;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11410;
 end   
18'd45203: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=43;
   mapp<=35;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12367;
 end   
18'd45204: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=68;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd45205: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=33;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd45206: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=95;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd45207: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=71;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd45208: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd45209: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd45210: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd45211: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd45212: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd45342: begin  
rid<=1;
end
18'd45343: begin  
end
18'd45344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd45345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd45346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd45347: begin  
rid<=0;
end
18'd45401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=12;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7479;
 end   
18'd45402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=93;
   mapp<=79;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4120;
 end   
18'd45403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd45404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd45405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd45542: begin  
rid<=1;
end
18'd45543: begin  
end
18'd45544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd45545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd45546: begin  
rid<=0;
end
18'd45601: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=6;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6600;
 end   
18'd45602: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=91;
   mapp<=58;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7886;
 end   
18'd45603: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=43;
   mapp<=26;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=7288;
 end   
18'd45604: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd45605: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=27;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd45606: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd45607: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd45608: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd45742: begin  
rid<=1;
end
18'd45743: begin  
end
18'd45744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd45745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd45746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd45747: begin  
rid<=0;
end
18'd45801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=67;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=20780;
 end   
18'd45802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=27;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=16443;
 end   
18'd45803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=5;
   mapp<=35;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=16358;
 end   
18'd45804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=46;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd45805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=86;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd45806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=89;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd45807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=40;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd45808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd45809: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd45810: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd45811: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd45812: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd45813: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20780;
 end   
18'd45814: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20780;
 end   
18'd45942: begin  
rid<=1;
end
18'd45943: begin  
end
18'd45944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd45945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd45946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd45947: begin  
rid<=0;
end
18'd46001: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=42;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4198;
 end   
18'd46002: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=0;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2680;
 end   
18'd46003: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=11;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd46004: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=25;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd46005: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=43;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd46006: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd46007: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd46008: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd46009: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd46142: begin  
rid<=1;
end
18'd46143: begin  
end
18'd46144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd46145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd46146: begin  
rid<=0;
end
18'd46201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=68;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1394;
 end   
18'd46202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=41;
   mapp<=4;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1353;
 end   
18'd46203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=35;
   mapp<=6;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1087;
 end   
18'd46204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=98;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=1678;
 end   
18'd46205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=25;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=605;
 end   
18'd46206: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=13;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd46207: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd46208: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd46209: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd46210: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd46342: begin  
rid<=1;
end
18'd46343: begin  
end
18'd46344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd46345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd46346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd46347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd46348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd46349: begin  
rid<=0;
end
18'd46401: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=46;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2622;
 end   
18'd46402: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=96;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=4426;
 end   
18'd46403: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=39;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=1814;
 end   
18'd46404: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=86;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=3986;
 end   
18'd46405: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=94;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=4364;
 end   
18'd46406: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd46542: begin  
rid<=1;
end
18'd46543: begin  
end
18'd46544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd46545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd46546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd46547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd46548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd46549: begin  
rid<=0;
end
18'd46601: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=90;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=18327;
 end   
18'd46602: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=73;
   mapp<=80;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=16372;
 end   
18'd46603: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=27;
   mapp<=55;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=16779;
 end   
18'd46604: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=13;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd46605: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=54;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd46606: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=96;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd46607: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=72;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd46608: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=50;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd46609: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd46610: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd46611: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd46612: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd46613: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18327;
 end   
18'd46614: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18327;
 end   
18'd46742: begin  
rid<=1;
end
18'd46743: begin  
end
18'd46744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd46745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd46746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd46747: begin  
rid<=0;
end
18'd46801: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=95;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9842;
 end   
18'd46802: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=3;
   mapp<=25;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7838;
 end   
18'd46803: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=94;
   mapp<=13;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=10788;
 end   
18'd46804: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=93;
   mapp<=24;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=10365;
 end   
18'd46805: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=67;
   mapp<=29;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=8902;
 end   
18'd46806: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=87;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=7788;
 end   
18'd46807: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=40;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=5994;
 end   
18'd46808: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=79;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd46809: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=41;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd46810: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=25;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd46811: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd46812: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd46813: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9842;
 end   
18'd46814: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9842;
 end   
18'd46815: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9842;
 end   
18'd46816: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9842;
 end   
18'd46942: begin  
rid<=1;
end
18'd46943: begin  
end
18'd46944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd46945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd46946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd46947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd46948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd46949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd46950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd46951: begin  
rid<=0;
end
18'd47001: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=11;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=20185;
 end   
18'd47002: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=25;
   mapp<=21;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=21487;
 end   
18'd47003: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=28;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd47004: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=78;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd47005: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=48;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd47006: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=50;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd47007: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=92;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd47008: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=44;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd47009: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=54;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd47010: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=23;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd47011: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=53;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd47012: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd47013: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20185;
 end   
18'd47014: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20185;
 end   
18'd47015: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20185;
 end   
18'd47016: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20185;
 end   
18'd47017: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20185;
 end   
18'd47018: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20185;
 end   
18'd47019: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20185;
 end   
18'd47020: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20185;
 end   
18'd47021: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20185;
 end   
18'd47142: begin  
rid<=1;
end
18'd47143: begin  
end
18'd47144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd47145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd47146: begin  
rid<=0;
end
18'd47201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=4;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5503;
 end   
18'd47202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=38;
   mapp<=26;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8850;
 end   
18'd47203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=71;
   mapp<=61;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5827;
 end   
18'd47204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=86;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=10155;
 end   
18'd47205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=5;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=6260;
 end   
18'd47206: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=99;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=7768;
 end   
18'd47207: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=56;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=7451;
 end   
18'd47208: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=28;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=6211;
 end   
18'd47209: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=67;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=5647;
 end   
18'd47210: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=51;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd47211: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=19;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd47212: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd47213: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5503;
 end   
18'd47214: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5503;
 end   
18'd47342: begin  
rid<=1;
end
18'd47343: begin  
end
18'd47344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd47345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd47346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd47347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd47348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd47349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd47350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd47351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd47352: begin  
check<=expctdoutput[8]-outcheck;
end
18'd47353: begin  
rid<=0;
end
18'd47401: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=12;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=18358;
 end   
18'd47402: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=67;
   mapp<=46;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=18255;
 end   
18'd47403: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=99;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd47404: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=44;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd47405: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=97;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd47406: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=1;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd47407: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd47408: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd47409: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd47410: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd47411: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd47542: begin  
rid<=1;
end
18'd47543: begin  
end
18'd47544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd47545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd47546: begin  
rid<=0;
end
18'd47601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=44;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16531;
 end   
18'd47602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=18;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13763;
 end   
18'd47603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=25;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd47604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=19;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd47605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=84;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd47606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=74;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd47607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd47608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd47609: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd47610: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd47611: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd47612: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd47613: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16531;
 end   
18'd47742: begin  
rid<=1;
end
18'd47743: begin  
end
18'd47744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd47745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd47746: begin  
rid<=0;
end
18'd47801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=14;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13288;
 end   
18'd47802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=63;
   mapp<=14;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11329;
 end   
18'd47803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=51;
   mapp<=95;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=18068;
 end   
18'd47804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=19;
   mapp<=3;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=10869;
 end   
18'd47805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=90;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd47806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=17;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd47807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=83;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd47808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=18;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd47809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=84;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd47810: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=52;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd47811: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd47812: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd47813: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13288;
 end   
18'd47814: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13288;
 end   
18'd47815: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13288;
 end   
18'd47816: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13288;
 end   
18'd47817: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13288;
 end   
18'd47942: begin  
rid<=1;
end
18'd47943: begin  
end
18'd47944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd47945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd47946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd47947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd47948: begin  
rid<=0;
end
18'd48001: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=37;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1776;
 end   
18'd48002: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=97;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4666;
 end   
18'd48003: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=24;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1172;
 end   
18'd48004: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=68;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=3294;
 end   
18'd48005: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=27;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=1336;
 end   
18'd48006: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=48;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=2354;
 end   
18'd48007: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=93;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=4524;
 end   
18'd48008: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=82;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=4006;
 end   
18'd48009: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd48142: begin  
rid<=1;
end
18'd48143: begin  
end
18'd48144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd48145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd48146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd48147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd48148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd48149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd48150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd48151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd48152: begin  
rid<=0;
end
18'd48201: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=77;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7161;
 end   
18'd48202: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=14;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1312;
 end   
18'd48203: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=4;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=392;
 end   
18'd48204: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=84;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=7842;
 end   
18'd48205: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=43;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=4039;
 end   
18'd48206: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd48342: begin  
rid<=1;
end
18'd48343: begin  
end
18'd48344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd48345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd48346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd48347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd48348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd48349: begin  
rid<=0;
end
18'd48401: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=92;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8556;
 end   
18'd48402: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=98;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9124;
 end   
18'd48403: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=90;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8390;
 end   
18'd48404: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=99;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=9237;
 end   
18'd48405: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=90;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=8410;
 end   
18'd48406: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd48542: begin  
rid<=1;
end
18'd48543: begin  
end
18'd48544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd48545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd48546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd48547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd48548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd48549: begin  
rid<=0;
end
18'd48601: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=14;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6088;
 end   
18'd48602: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=73;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd48603: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd48604: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd48742: begin  
rid<=1;
end
18'd48743: begin  
end
18'd48744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd48745: begin  
rid<=0;
end
18'd48801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=38;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2833;
 end   
18'd48802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=11;
   mapp<=33;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2441;
 end   
18'd48803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=52;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd48804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd48805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd48942: begin  
rid<=1;
end
18'd48943: begin  
end
18'd48944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd48945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd48946: begin  
rid<=0;
end
18'd49001: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=68;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13687;
 end   
18'd49002: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=21;
   mapp<=88;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13595;
 end   
18'd49003: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=58;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd49004: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=57;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd49005: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=47;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd49006: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=82;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd49007: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=38;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd49008: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=22;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd49009: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd49010: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd49011: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd49012: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd49013: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13687;
 end   
18'd49014: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13687;
 end   
18'd49015: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13687;
 end   
18'd49142: begin  
rid<=1;
end
18'd49143: begin  
end
18'd49144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd49145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd49146: begin  
rid<=0;
end
18'd49201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=45;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6097;
 end   
18'd49202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=51;
   mapp<=89;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3371;
 end   
18'd49203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=23;
   mapp<=56;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=4560;
 end   
18'd49204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=18;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd49205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=50;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd49206: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd49207: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd49208: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd49342: begin  
rid<=1;
end
18'd49343: begin  
end
18'd49344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd49345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd49346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd49347: begin  
rid<=0;
end
18'd49401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=41;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3731;
 end   
18'd49402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=6;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=256;
 end   
18'd49403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=10;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=430;
 end   
18'd49404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=13;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=563;
 end   
18'd49405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=51;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=2131;
 end   
18'd49406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=80;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=3330;
 end   
18'd49407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=44;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=1864;
 end   
18'd49408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=43;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=1833;
 end   
18'd49409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd49542: begin  
rid<=1;
end
18'd49543: begin  
end
18'd49544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd49545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd49546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd49547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd49548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd49549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd49550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd49551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd49552: begin  
rid<=0;
end
18'd49601: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=27;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6259;
 end   
18'd49602: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=24;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd49603: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=4;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd49604: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=56;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd49605: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd49606: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd49607: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd49608: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd49742: begin  
rid<=1;
end
18'd49743: begin  
end
18'd49744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd49745: begin  
rid<=0;
end
18'd49801: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=98;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5548;
 end   
18'd49802: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=79;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7000;
 end   
18'd49803: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=86;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=13820;
 end   
18'd49804: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd49805: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd49806: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd49942: begin  
rid<=1;
end
18'd49943: begin  
end
18'd49944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd49945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd49946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd49947: begin  
rid<=0;
end
18'd50001: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=96;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12116;
 end   
18'd50002: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=50;
   mapp<=90;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=15805;
 end   
18'd50003: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=12;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd50004: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=22;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd50005: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=29;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd50006: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd50007: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd50008: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd50009: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd50010: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd50011: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd50142: begin  
rid<=1;
end
18'd50143: begin  
end
18'd50144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd50145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd50146: begin  
rid<=0;
end
18'd50201: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=51;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=20825;
 end   
18'd50202: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=97;
   mapp<=53;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=24357;
 end   
18'd50203: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=51;
   mapp<=76;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=20122;
 end   
18'd50204: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=1;
   mapp<=70;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=16262;
 end   
18'd50205: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=35;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd50206: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=93;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd50207: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=72;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd50208: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd50209: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd50210: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd50211: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd50212: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd50213: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20825;
 end   
18'd50214: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20825;
 end   
18'd50215: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20825;
 end   
18'd50342: begin  
rid<=1;
end
18'd50343: begin  
end
18'd50344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd50345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd50346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd50347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd50348: begin  
rid<=0;
end
18'd50401: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=2;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15305;
 end   
18'd50402: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=58;
   mapp<=38;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=14826;
 end   
18'd50403: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=88;
   mapp<=96;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9758;
 end   
18'd50404: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=21;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd50405: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=86;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd50406: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd50407: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd50408: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd50409: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd50410: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd50411: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd50412: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd50542: begin  
rid<=1;
end
18'd50543: begin  
end
18'd50544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd50545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd50546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd50547: begin  
rid<=0;
end
18'd50601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=62;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1736;
 end   
18'd50602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=79;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=4908;
 end   
18'd50603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=47;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=2934;
 end   
18'd50604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=49;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=3068;
 end   
18'd50605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=80;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=5000;
 end   
18'd50606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=45;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=2840;
 end   
18'd50607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=28;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=1796;
 end   
18'd50608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd50742: begin  
rid<=1;
end
18'd50743: begin  
end
18'd50744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd50745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd50746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd50747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd50748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd50749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd50750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd50751: begin  
rid<=0;
end
18'd50801: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=56;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4312;
 end   
18'd50802: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=91;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=5106;
 end   
18'd50803: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=47;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=2652;
 end   
18'd50804: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=85;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=4790;
 end   
18'd50805: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=31;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=1776;
 end   
18'd50806: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=6;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=386;
 end   
18'd50807: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=84;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=4764;
 end   
18'd50808: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=54;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=3094;
 end   
18'd50809: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=69;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=3944;
 end   
18'd50810: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=9;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[9]<=594;
 end   
18'd50811: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd50942: begin  
rid<=1;
end
18'd50943: begin  
end
18'd50944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd50945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd50946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd50947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd50948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd50949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd50950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd50951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd50952: begin  
check<=expctdoutput[8]-outcheck;
end
18'd50953: begin  
check<=expctdoutput[9]-outcheck;
end
18'd50954: begin  
rid<=0;
end
18'd51001: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=35;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13088;
 end   
18'd51002: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=90;
   mapp<=16;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10517;
 end   
18'd51003: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=77;
   mapp<=60;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=14451;
 end   
18'd51004: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=49;
   mapp<=97;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=16991;
 end   
18'd51005: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=5;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd51006: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=86;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd51007: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd51008: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd51009: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd51010: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd51011: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd51142: begin  
rid<=1;
end
18'd51143: begin  
end
18'd51144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd51145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd51146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd51147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd51148: begin  
rid<=0;
end
18'd51201: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=88;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=22183;
 end   
18'd51202: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=15;
   mapp<=30;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=21006;
 end   
18'd51203: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=8;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd51204: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=10;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd51205: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=40;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd51206: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=99;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd51207: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=97;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd51208: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=7;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd51209: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=54;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd51210: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=4;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd51211: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd51212: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd51213: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22183;
 end   
18'd51214: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22183;
 end   
18'd51215: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22183;
 end   
18'd51216: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22183;
 end   
18'd51217: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22183;
 end   
18'd51218: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22183;
 end   
18'd51219: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22183;
 end   
18'd51342: begin  
rid<=1;
end
18'd51343: begin  
end
18'd51344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd51345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd51346: begin  
rid<=0;
end
18'd51401: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6967;
 end   
18'd51402: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=64;
   mapp<=92;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1838;
 end   
18'd51403: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=83;
   mapp<=13;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=7594;
 end   
18'd51404: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=12;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=12167;
 end   
18'd51405: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=82;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=9585;
 end   
18'd51406: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=83;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=5721;
 end   
18'd51407: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=51;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=4987;
 end   
18'd51408: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=29;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=5177;
 end   
18'd51409: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd51410: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd51411: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd51412: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd51413: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6967;
 end   
18'd51542: begin  
rid<=1;
end
18'd51543: begin  
end
18'd51544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd51545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd51546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd51547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd51548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd51549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd51550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd51551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd51552: begin  
rid<=0;
end
18'd51601: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=56;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10703;
 end   
18'd51602: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=92;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8978;
 end   
18'd51603: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=40;
   mapp<=8;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8739;
 end   
18'd51604: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=87;
   mapp<=41;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=14058;
 end   
18'd51605: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=32;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=17209;
 end   
18'd51606: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=37;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=13897;
 end   
18'd51607: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=84;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=19915;
 end   
18'd51608: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=99;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=15687;
 end   
18'd51609: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd51610: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd51611: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd51612: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd51613: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10703;
 end   
18'd51614: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10703;
 end   
18'd51615: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10703;
 end   
18'd51742: begin  
rid<=1;
end
18'd51743: begin  
end
18'd51744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd51745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd51746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd51747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd51748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd51749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd51750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd51751: begin  
check<=expctdoutput[7]-outcheck;
end
18'd51752: begin  
rid<=0;
end
18'd51801: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=33;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=18241;
 end   
18'd51802: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=78;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=17865;
 end   
18'd51803: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=86;
   mapp<=63;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=18525;
 end   
18'd51804: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=24;
   mapp<=15;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=21620;
 end   
18'd51805: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=34;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd51806: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=75;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd51807: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd51808: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd51809: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd51810: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd51811: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd51812: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd51813: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18241;
 end   
18'd51814: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18241;
 end   
18'd51815: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18241;
 end   
18'd51942: begin  
rid<=1;
end
18'd51943: begin  
end
18'd51944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd51945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd51946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd51947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd51948: begin  
rid<=0;
end
18'd52001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=55;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4620;
 end   
18'd52002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=24;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=1330;
 end   
18'd52003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=92;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=5080;
 end   
18'd52004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=4;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=250;
 end   
18'd52005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=22;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=1250;
 end   
18'd52006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd52142: begin  
rid<=1;
end
18'd52143: begin  
end
18'd52144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd52145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd52146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd52147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd52148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd52149: begin  
rid<=0;
end
18'd52201: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=97;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7081;
 end   
18'd52202: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=84;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=8158;
 end   
18'd52203: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=60;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=5840;
 end   
18'd52204: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=22;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=2164;
 end   
18'd52205: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=53;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=5181;
 end   
18'd52206: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd52342: begin  
rid<=1;
end
18'd52343: begin  
end
18'd52344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd52345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd52346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd52347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd52348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd52349: begin  
rid<=0;
end
18'd52401: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=90;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15571;
 end   
18'd52402: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=98;
   mapp<=17;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13054;
 end   
18'd52403: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=85;
   mapp<=6;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=20346;
 end   
18'd52404: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=47;
   mapp<=31;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=28339;
 end   
18'd52405: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=84;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd52406: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=92;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd52407: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd52408: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd52409: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd52410: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd52411: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd52412: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd52413: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15571;
 end   
18'd52414: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15571;
 end   
18'd52415: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15571;
 end   
18'd52542: begin  
rid<=1;
end
18'd52543: begin  
end
18'd52544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd52545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd52546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd52547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd52548: begin  
rid<=0;
end
18'd52601: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=28;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7350;
 end   
18'd52602: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=95;
   mapp<=28;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8069;
 end   
18'd52603: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=42;
   mapp<=38;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6408;
 end   
18'd52604: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=37;
   mapp<=42;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=7005;
 end   
18'd52605: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=6;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=8166;
 end   
18'd52606: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=67;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=8963;
 end   
18'd52607: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=53;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=7701;
 end   
18'd52608: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=93;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd52609: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=5;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd52610: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=46;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd52611: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd52612: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd52613: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7350;
 end   
18'd52614: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7350;
 end   
18'd52742: begin  
rid<=1;
end
18'd52743: begin  
end
18'd52744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd52745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd52746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd52747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd52748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd52749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd52750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd52751: begin  
rid<=0;
end
18'd52801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=39;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2496;
 end   
18'd52802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=6;
   mapp<=65;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=919;
 end   
18'd52803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=9;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6486;
 end   
18'd52804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=92;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=11433;
 end   
18'd52805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=99;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=10261;
 end   
18'd52806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=75;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=6440;
 end   
18'd52807: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=36;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=5969;
 end   
18'd52808: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=61;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=6419;
 end   
18'd52809: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=47;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=3788;
 end   
18'd52810: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=18;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd52811: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd52812: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd52942: begin  
rid<=1;
end
18'd52943: begin  
end
18'd52944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd52945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd52946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd52947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd52948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd52949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd52950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd52951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd52952: begin  
check<=expctdoutput[8]-outcheck;
end
18'd52953: begin  
rid<=0;
end
18'd53001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=44;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=21869;
 end   
18'd53002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=36;
   mapp<=96;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=23211;
 end   
18'd53003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=37;
   mapp<=9;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=20539;
 end   
18'd53004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=16;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd53005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=93;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd53006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=49;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd53007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=71;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd53008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=44;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd53009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=77;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd53010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd53011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd53012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd53013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21869;
 end   
18'd53014: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21869;
 end   
18'd53015: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21869;
 end   
18'd53016: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21869;
 end   
18'd53017: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21869;
 end   
18'd53018: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21869;
 end   
18'd53019: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21869;
 end   
18'd53020: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21869;
 end   
18'd53142: begin  
rid<=1;
end
18'd53143: begin  
end
18'd53144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd53145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd53146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd53147: begin  
rid<=0;
end
18'd53201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=18;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7550;
 end   
18'd53202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=68;
   mapp<=85;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7365;
 end   
18'd53203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=6;
   mapp<=25;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=3225;
 end   
18'd53204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=29;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=4345;
 end   
18'd53205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=8;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=4870;
 end   
18'd53206: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=41;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=6765;
 end   
18'd53207: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=25;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=7370;
 end   
18'd53208: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=36;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=10510;
 end   
18'd53209: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=80;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd53210: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd53211: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd53212: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd53213: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7550;
 end   
18'd53342: begin  
rid<=1;
end
18'd53343: begin  
end
18'd53344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd53345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd53346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd53347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd53348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd53349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd53350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd53351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd53352: begin  
rid<=0;
end
18'd53401: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=28;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1316;
 end   
18'd53402: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=36;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1702;
 end   
18'd53403: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=4;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=208;
 end   
18'd53404: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=30;
 end   
18'd53405: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=23;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=1121;
 end   
18'd53406: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=64;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=3058;
 end   
18'd53407: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=11;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=577;
 end   
18'd53408: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd53542: begin  
rid<=1;
end
18'd53543: begin  
end
18'd53544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd53545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd53546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd53547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd53548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd53549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd53550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd53551: begin  
rid<=0;
end
18'd53601: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=41;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8944;
 end   
18'd53602: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=70;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4421;
 end   
18'd53603: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=45;
   mapp<=66;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6506;
 end   
18'd53604: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=6;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=11054;
 end   
18'd53605: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=88;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=5502;
 end   
18'd53606: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=56;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=5211;
 end   
18'd53607: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=7;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=9328;
 end   
18'd53608: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=66;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd53609: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=57;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd53610: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd53611: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd53612: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd53742: begin  
rid<=1;
end
18'd53743: begin  
end
18'd53744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd53745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd53746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd53747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd53748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd53749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd53750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd53751: begin  
rid<=0;
end
18'd53801: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=90;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=19965;
 end   
18'd53802: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=67;
   mapp<=55;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=18873;
 end   
18'd53803: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=7;
   mapp<=91;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=18611;
 end   
18'd53804: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=34;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd53805: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=46;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd53806: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=62;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd53807: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=2;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd53808: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=39;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd53809: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=26;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd53810: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=95;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd53811: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd53812: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd53813: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19965;
 end   
18'd53814: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19965;
 end   
18'd53815: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19965;
 end   
18'd53816: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19965;
 end   
18'd53817: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19965;
 end   
18'd53818: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19965;
 end   
18'd53942: begin  
rid<=1;
end
18'd53943: begin  
end
18'd53944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd53945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd53946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd53947: begin  
rid<=0;
end
18'd54001: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=76;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=21687;
 end   
18'd54002: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=64;
   mapp<=86;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=21291;
 end   
18'd54003: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=57;
   mapp<=79;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=18671;
 end   
18'd54004: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=70;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd54005: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=38;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd54006: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=12;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd54007: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=44;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd54008: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=61;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd54009: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=80;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd54010: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd54011: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd54012: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd54013: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21687;
 end   
18'd54014: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21687;
 end   
18'd54015: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21687;
 end   
18'd54016: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21687;
 end   
18'd54017: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21687;
 end   
18'd54018: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21687;
 end   
18'd54142: begin  
rid<=1;
end
18'd54143: begin  
end
18'd54144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd54145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd54146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd54147: begin  
rid<=0;
end
18'd54201: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=7;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=17037;
 end   
18'd54202: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=84;
   mapp<=47;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=19690;
 end   
18'd54203: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=47;
   mapp<=39;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=18741;
 end   
18'd54204: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=77;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd54205: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=75;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd54206: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=13;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd54207: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=9;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd54208: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=71;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd54209: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=42;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd54210: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=39;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd54211: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=36;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd54212: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd54213: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17037;
 end   
18'd54214: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17037;
 end   
18'd54215: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17037;
 end   
18'd54216: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17037;
 end   
18'd54217: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17037;
 end   
18'd54218: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17037;
 end   
18'd54219: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17037;
 end   
18'd54220: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17037;
 end   
18'd54342: begin  
rid<=1;
end
18'd54343: begin  
end
18'd54344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd54345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd54346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd54347: begin  
rid<=0;
end
18'd54401: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=98;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13625;
 end   
18'd54402: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=2;
   mapp<=29;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9940;
 end   
18'd54403: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=5;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd54404: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=38;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd54405: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=32;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd54406: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=65;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd54407: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=16;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd54408: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=81;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd54409: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd54410: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd54411: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd54412: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd54413: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13625;
 end   
18'd54414: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13625;
 end   
18'd54415: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13625;
 end   
18'd54542: begin  
rid<=1;
end
18'd54543: begin  
end
18'd54544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd54545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd54546: begin  
rid<=0;
end
18'd54601: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=40;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4918;
 end   
18'd54602: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=16;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd54603: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=88;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd54604: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=19;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd54605: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd54606: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd54607: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd54608: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd54742: begin  
rid<=1;
end
18'd54743: begin  
end
18'd54744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd54745: begin  
rid<=0;
end
18'd54801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=71;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8422;
 end   
18'd54802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=83;
   mapp<=51;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8171;
 end   
18'd54803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=64;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd54804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd54805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd54942: begin  
rid<=1;
end
18'd54943: begin  
end
18'd54944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd54945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd54946: begin  
rid<=0;
end
18'd55001: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=59;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4956;
 end   
18'd55002: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=1;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=94;
 end   
18'd55003: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=74;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6236;
 end   
18'd55004: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=33;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=2802;
 end   
18'd55005: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=59;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=4996;
 end   
18'd55006: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=14;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=1226;
 end   
18'd55007: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=49;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=4176;
 end   
18'd55008: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=95;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=8050;
 end   
18'd55009: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=22;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=1928;
 end   
18'd55010: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=41;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[9]<=3534;
 end   
18'd55011: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd55142: begin  
rid<=1;
end
18'd55143: begin  
end
18'd55144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd55145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd55146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd55147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd55148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd55149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd55150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd55151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd55152: begin  
check<=expctdoutput[8]-outcheck;
end
18'd55153: begin  
check<=expctdoutput[9]-outcheck;
end
18'd55154: begin  
rid<=0;
end
18'd55201: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=65;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3380;
 end   
18'd55202: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=91;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4742;
 end   
18'd55203: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=38;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1996;
 end   
18'd55204: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=10;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=550;
 end   
18'd55205: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=67;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=3524;
 end   
18'd55206: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=55;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=2910;
 end   
18'd55207: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=87;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=4584;
 end   
18'd55208: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=24;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=1318;
 end   
18'd55209: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=22;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=1224;
 end   
18'd55210: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=39;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[9]<=2118;
 end   
18'd55211: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=41;
   mapp<=0;
   pp<=100;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[10]<=2232;
 end   
18'd55212: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd55342: begin  
rid<=1;
end
18'd55343: begin  
end
18'd55344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd55345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd55346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd55347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd55348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd55349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd55350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd55351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd55352: begin  
check<=expctdoutput[8]-outcheck;
end
18'd55353: begin  
check<=expctdoutput[9]-outcheck;
end
18'd55354: begin  
check<=expctdoutput[10]-outcheck;
end
18'd55355: begin  
rid<=0;
end
18'd55401: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=74;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14365;
 end   
18'd55402: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=76;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=12475;
 end   
18'd55403: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=37;
   mapp<=41;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9667;
 end   
18'd55404: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=33;
   mapp<=72;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=8101;
 end   
18'd55405: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=41;
   mapp<=68;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=11344;
 end   
18'd55406: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=45;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd55407: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=18;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd55408: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=15;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd55409: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=74;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd55410: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd55411: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd55412: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd55413: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14365;
 end   
18'd55414: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14365;
 end   
18'd55542: begin  
rid<=1;
end
18'd55543: begin  
end
18'd55544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd55545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd55546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd55547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd55548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd55549: begin  
rid<=0;
end
18'd55601: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=81;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8232;
 end   
18'd55602: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=44;
   mapp<=24;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5678;
 end   
18'd55603: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=40;
   mapp<=66;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9412;
 end   
18'd55604: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=34;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=9254;
 end   
18'd55605: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=96;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=9022;
 end   
18'd55606: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=76;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=5284;
 end   
18'd55607: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=27;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=2880;
 end   
18'd55608: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=5;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=6788;
 end   
18'd55609: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=18;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=5978;
 end   
18'd55610: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=91;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd55611: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=41;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd55612: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd55613: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8232;
 end   
18'd55614: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8232;
 end   
18'd55742: begin  
rid<=1;
end
18'd55743: begin  
end
18'd55744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd55745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd55746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd55747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd55748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd55749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd55750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd55751: begin  
check<=expctdoutput[7]-outcheck;
end
18'd55752: begin  
check<=expctdoutput[8]-outcheck;
end
18'd55753: begin  
rid<=0;
end
18'd55801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=0;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1003;
 end   
18'd55802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=17;
   mapp<=59;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2161;
 end   
18'd55803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=16;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=3693;
 end   
18'd55804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=43;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=4499;
 end   
18'd55805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=24;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=5520;
 end   
18'd55806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=64;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=4889;
 end   
18'd55807: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=5;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=3778;
 end   
18'd55808: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=57;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=4235;
 end   
18'd55809: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=2;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=4116;
 end   
18'd55810: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=66;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[9]<=9201;
 end   
18'd55811: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=75;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd55812: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd55813: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=1003;
 end   
18'd55942: begin  
rid<=1;
end
18'd55943: begin  
end
18'd55944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd55945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd55946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd55947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd55948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd55949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd55950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd55951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd55952: begin  
check<=expctdoutput[8]-outcheck;
end
18'd55953: begin  
check<=expctdoutput[9]-outcheck;
end
18'd55954: begin  
rid<=0;
end
18'd56001: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=52;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6003;
 end   
18'd56002: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=1;
   mapp<=46;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3932;
 end   
18'd56003: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=26;
   mapp<=45;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8699;
 end   
18'd56004: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=53;
   mapp<=3;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=10966;
 end   
18'd56005: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=84;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=12035;
 end   
18'd56006: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=49;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=7074;
 end   
18'd56007: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=50;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=6885;
 end   
18'd56008: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=5;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=3966;
 end   
18'd56009: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=46;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd56010: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=25;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd56011: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd56012: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd56013: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6003;
 end   
18'd56014: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6003;
 end   
18'd56015: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6003;
 end   
18'd56142: begin  
rid<=1;
end
18'd56143: begin  
end
18'd56144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd56145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd56146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd56147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd56148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd56149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd56150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd56151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd56152: begin  
rid<=0;
end
18'd56201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=96;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16742;
 end   
18'd56202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=10;
   mapp<=23;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8432;
 end   
18'd56203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=76;
   mapp<=32;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=15844;
 end   
18'd56204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=92;
   mapp<=56;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=17936;
 end   
18'd56205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=50;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=12712;
 end   
18'd56206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=90;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=15069;
 end   
18'd56207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=95;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=12531;
 end   
18'd56208: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=52;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=8552;
 end   
18'd56209: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=50;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd56210: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=15;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd56211: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=36;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd56212: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd56213: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16742;
 end   
18'd56214: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16742;
 end   
18'd56215: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16742;
 end   
18'd56342: begin  
rid<=1;
end
18'd56343: begin  
end
18'd56344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd56345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd56346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd56347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd56348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd56349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd56350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd56351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd56352: begin  
rid<=0;
end
18'd56401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=50;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6782;
 end   
18'd56402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=82;
   mapp<=29;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8296;
 end   
18'd56403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=6;
   mapp<=34;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=4424;
 end   
18'd56404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=36;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=8550;
 end   
18'd56405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=84;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=10284;
 end   
18'd56406: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=90;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=10891;
 end   
18'd56407: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=17;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=6110;
 end   
18'd56408: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=82;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=9416;
 end   
18'd56409: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=66;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd56410: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd56411: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd56412: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd56413: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6782;
 end   
18'd56542: begin  
rid<=1;
end
18'd56543: begin  
end
18'd56544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd56545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd56546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd56547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd56548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd56549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd56550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd56551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd56552: begin  
rid<=0;
end
18'd56601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=95;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=28486;
 end   
18'd56602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=80;
   mapp<=10;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=24847;
 end   
18'd56603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=38;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd56604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=67;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd56605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=20;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd56606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=45;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd56607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=83;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd56608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=65;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd56609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=96;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd56610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=33;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd56611: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd56612: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd56613: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28486;
 end   
18'd56614: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28486;
 end   
18'd56615: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28486;
 end   
18'd56616: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28486;
 end   
18'd56617: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28486;
 end   
18'd56618: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28486;
 end   
18'd56619: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28486;
 end   
18'd56742: begin  
rid<=1;
end
18'd56743: begin  
end
18'd56744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd56745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd56746: begin  
rid<=0;
end
18'd56801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=13;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10710;
 end   
18'd56802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=39;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9968;
 end   
18'd56803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=52;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd56804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=45;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd56805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=61;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd56806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=51;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd56807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd56808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd56809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd56810: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd56811: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd56812: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd56813: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10710;
 end   
18'd56942: begin  
rid<=1;
end
18'd56943: begin  
end
18'd56944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd56945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd56946: begin  
rid<=0;
end
18'd57001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=11;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=143;
 end   
18'd57002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=7;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=87;
 end   
18'd57003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=54;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=614;
 end   
18'd57004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=76;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=866;
 end   
18'd57005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=17;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=227;
 end   
18'd57006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd57142: begin  
rid<=1;
end
18'd57143: begin  
end
18'd57144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd57145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd57146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd57147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd57148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd57149: begin  
rid<=0;
end
18'd57201: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=64;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=27501;
 end   
18'd57202: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=62;
   mapp<=31;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=29957;
 end   
18'd57203: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=10;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd57204: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=46;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd57205: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=65;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd57206: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=80;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd57207: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=65;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd57208: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=46;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd57209: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=40;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd57210: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=97;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd57211: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd57212: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd57213: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=27501;
 end   
18'd57214: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=27501;
 end   
18'd57215: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=27501;
 end   
18'd57216: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=27501;
 end   
18'd57217: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=27501;
 end   
18'd57218: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=27501;
 end   
18'd57219: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=27501;
 end   
18'd57342: begin  
rid<=1;
end
18'd57343: begin  
end
18'd57344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd57345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd57346: begin  
rid<=0;
end
18'd57401: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=70;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7840;
 end   
18'd57402: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=15;
   mapp<=84;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1420;
 end   
18'd57403: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=524;
 end   
18'd57404: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=6;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=1098;
 end   
18'd57405: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=6;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=772;
 end   
18'd57406: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=2;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=8302;
 end   
18'd57407: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=96;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=11856;
 end   
18'd57408: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=33;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=4096;
 end   
18'd57409: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=11;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=6742;
 end   
18'd57410: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=67;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[9]<=7648;
 end   
18'd57411: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=15;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd57412: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd57413: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7840;
 end   
18'd57542: begin  
rid<=1;
end
18'd57543: begin  
end
18'd57544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd57545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd57546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd57547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd57548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd57549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd57550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd57551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd57552: begin  
check<=expctdoutput[8]-outcheck;
end
18'd57553: begin  
check<=expctdoutput[9]-outcheck;
end
18'd57554: begin  
rid<=0;
end
18'd57601: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=19;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4818;
 end   
18'd57602: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=79;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8500;
 end   
18'd57603: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd57604: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd57605: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd57742: begin  
rid<=1;
end
18'd57743: begin  
end
18'd57744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd57745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd57746: begin  
rid<=0;
end
18'd57801: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=99;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11723;
 end   
18'd57802: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=20;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10833;
 end   
18'd57803: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=20;
   mapp<=9;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=3371;
 end   
18'd57804: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=52;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=7758;
 end   
18'd57805: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=71;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=8669;
 end   
18'd57806: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=58;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=7412;
 end   
18'd57807: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=22;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=5358;
 end   
18'd57808: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=59;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=9831;
 end   
18'd57809: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd57810: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd57811: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd57812: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd57813: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11723;
 end   
18'd57942: begin  
rid<=1;
end
18'd57943: begin  
end
18'd57944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd57945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd57946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd57947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd57948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd57949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd57950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd57951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd57952: begin  
rid<=0;
end
18'd58001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=99;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1188;
 end   
18'd58002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=15;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=1495;
 end   
18'd58003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=53;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=5267;
 end   
18'd58004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=85;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=8445;
 end   
18'd58005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=41;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=4099;
 end   
18'd58006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd58142: begin  
rid<=1;
end
18'd58143: begin  
end
18'd58144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd58145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd58146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd58147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd58148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd58149: begin  
rid<=0;
end
18'd58201: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=6;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16381;
 end   
18'd58202: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=49;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd58203: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=75;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd58204: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=26;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd58205: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=24;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd58206: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=7;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd58207: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=74;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd58208: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd58209: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd58210: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd58211: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd58212: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd58213: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16381;
 end   
18'd58214: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16381;
 end   
18'd58342: begin  
rid<=1;
end
18'd58343: begin  
end
18'd58344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd58345: begin  
rid<=0;
end
18'd58401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=14;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8357;
 end   
18'd58402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=49;
   mapp<=45;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8402;
 end   
18'd58403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=68;
   mapp<=81;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5425;
 end   
18'd58404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=38;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=9626;
 end   
18'd58405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=7;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=4871;
 end   
18'd58406: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=93;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=4913;
 end   
18'd58407: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=4;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=8326;
 end   
18'd58408: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=5;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=6042;
 end   
18'd58409: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=97;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd58410: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=17;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd58411: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd58412: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd58413: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8357;
 end   
18'd58542: begin  
rid<=1;
end
18'd58543: begin  
end
18'd58544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd58545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd58546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd58547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd58548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd58549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd58550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd58551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd58552: begin  
rid<=0;
end
18'd58601: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=33;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14708;
 end   
18'd58602: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=54;
   mapp<=33;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=16366;
 end   
18'd58603: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=30;
   mapp<=97;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=16673;
 end   
18'd58604: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=52;
   mapp<=79;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=22503;
 end   
18'd58605: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=4;
   mapp<=36;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=22789;
 end   
18'd58606: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=79;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd58607: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd58608: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd58609: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=54;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd58610: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=72;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd58611: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd58612: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd58613: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14708;
 end   
18'd58614: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14708;
 end   
18'd58615: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14708;
 end   
18'd58616: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14708;
 end   
18'd58742: begin  
rid<=1;
end
18'd58743: begin  
end
18'd58744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd58745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd58746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd58747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd58748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd58749: begin  
rid<=0;
end
18'd58801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=31;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7345;
 end   
18'd58802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=80;
   mapp<=86;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7660;
 end   
18'd58803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=75;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6305;
 end   
18'd58804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=60;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=2134;
 end   
18'd58805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=14;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd58806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd58807: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd58942: begin  
rid<=1;
end
18'd58943: begin  
end
18'd58944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd58945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd58946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd58947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd58948: begin  
rid<=0;
end
18'd59001: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=31;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10454;
 end   
18'd59002: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=61;
   mapp<=38;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10424;
 end   
18'd59003: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=19;
   mapp<=81;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=7654;
 end   
18'd59004: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=81;
   mapp<=47;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=10061;
 end   
18'd59005: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd59006: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd59007: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd59008: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd59009: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd59010: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd59011: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd59142: begin  
rid<=1;
end
18'd59143: begin  
end
18'd59144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd59145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd59146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd59147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd59148: begin  
rid<=0;
end
18'd59201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=2;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1950;
 end   
18'd59202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=28;
   mapp<=63;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3545;
 end   
18'd59203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=21;
   mapp<=2;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=7800;
 end   
18'd59204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=98;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=10137;
 end   
18'd59205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=47;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=6271;
 end   
18'd59206: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=45;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=3712;
 end   
18'd59207: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=6;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd59208: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=22;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd59209: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd59210: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd59211: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd59342: begin  
rid<=1;
end
18'd59343: begin  
end
18'd59344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd59345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd59346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd59347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd59348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd59349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd59350: begin  
rid<=0;
end
18'd59401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=37;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=24033;
 end   
18'd59402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=53;
   mapp<=44;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=21784;
 end   
18'd59403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=68;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd59404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=30;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd59405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=55;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd59406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=66;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd59407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=58;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd59408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=12;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd59409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=56;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd59410: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd59411: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd59412: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd59413: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24033;
 end   
18'd59414: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24033;
 end   
18'd59415: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24033;
 end   
18'd59416: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24033;
 end   
18'd59417: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24033;
 end   
18'd59542: begin  
rid<=1;
end
18'd59543: begin  
end
18'd59544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd59545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd59546: begin  
rid<=0;
end
18'd59601: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=50;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7800;
 end   
18'd59602: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=75;
   mapp<=76;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4260;
 end   
18'd59603: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=6;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=470;
 end   
18'd59604: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=2;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=6430;
 end   
18'd59605: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=84;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=5965;
 end   
18'd59606: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=23;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=6450;
 end   
18'd59607: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=70;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=4460;
 end   
18'd59608: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd59609: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd59610: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd59742: begin  
rid<=1;
end
18'd59743: begin  
end
18'd59744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd59745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd59746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd59747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd59748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd59749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd59750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd59751: begin  
rid<=0;
end
18'd59801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=92;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=27986;
 end   
18'd59802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=48;
   mapp<=88;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=22309;
 end   
18'd59803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=84;
   mapp<=20;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=23015;
 end   
18'd59804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=45;
   mapp<=1;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=23840;
 end   
18'd59805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=87;
   mapp<=83;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=26534;
 end   
18'd59806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=62;
   mapp<=98;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=18404;
 end   
18'd59807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=43;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd59808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=58;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd59809: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=59;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd59810: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=71;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd59811: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd59812: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd59813: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=27986;
 end   
18'd59814: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=27986;
 end   
18'd59815: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=27986;
 end   
18'd59816: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=27986;
 end   
18'd59817: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=27986;
 end   
18'd59942: begin  
rid<=1;
end
18'd59943: begin  
end
18'd59944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd59945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd59946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd59947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd59948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd59949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd59950: begin  
rid<=0;
end
18'd60001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=46;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=25978;
 end   
18'd60002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=69;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=20325;
 end   
18'd60003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=75;
   mapp<=88;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=23081;
 end   
18'd60004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=17;
   mapp<=15;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=18107;
 end   
18'd60005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=87;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd60006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=20;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd60007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=30;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd60008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=42;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd60009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd60010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd60011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd60012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd60013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25978;
 end   
18'd60014: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25978;
 end   
18'd60015: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25978;
 end   
18'd60016: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25978;
 end   
18'd60017: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25978;
 end   
18'd60018: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25978;
 end   
18'd60019: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25978;
 end   
18'd60142: begin  
rid<=1;
end
18'd60143: begin  
end
18'd60144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd60145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd60146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd60147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd60148: begin  
rid<=0;
end
18'd60201: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=13;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=27867;
 end   
18'd60202: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=35;
   mapp<=80;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=28564;
 end   
18'd60203: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=35;
   mapp<=73;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=22819;
 end   
18'd60204: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=83;
   mapp<=77;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=20143;
 end   
18'd60205: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=86;
   mapp<=86;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=20248;
 end   
18'd60206: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=96;
   mapp<=81;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=23537;
 end   
18'd60207: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd60208: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd60209: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd60210: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd60211: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd60212: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd60213: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=27867;
 end   
18'd60214: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=27867;
 end   
18'd60215: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=27867;
 end   
18'd60216: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=27867;
 end   
18'd60217: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=27867;
 end   
18'd60342: begin  
rid<=1;
end
18'd60343: begin  
end
18'd60344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd60345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd60346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd60347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd60348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd60349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd60350: begin  
rid<=0;
end
18'd60401: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=60;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4842;
 end   
18'd60402: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=82;
   mapp<=21;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5030;
 end   
18'd60403: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=36;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=3740;
 end   
18'd60404: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=88;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=5005;
 end   
18'd60405: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=19;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=1784;
 end   
18'd60406: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=36;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=3854;
 end   
18'd60407: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=92;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd60408: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd60409: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd60542: begin  
rid<=1;
end
18'd60543: begin  
end
18'd60544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd60545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd60546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd60547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd60548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd60549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd60550: begin  
rid<=0;
end
18'd60601: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=21;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12839;
 end   
18'd60602: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=2;
   mapp<=96;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11750;
 end   
18'd60603: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=45;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd60604: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=2;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd60605: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=64;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd60606: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=39;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd60607: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=72;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd60608: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd60609: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd60610: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd60611: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd60612: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd60613: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12839;
 end   
18'd60742: begin  
rid<=1;
end
18'd60743: begin  
end
18'd60744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd60745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd60746: begin  
rid<=0;
end
18'd60801: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=80;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12261;
 end   
18'd60802: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=98;
   mapp<=54;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10424;
 end   
18'd60803: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=91;
   mapp<=59;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5670;
 end   
18'd60804: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=60;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=7139;
 end   
18'd60805: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=10;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd60806: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=91;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd60807: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd60808: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd60809: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd60942: begin  
rid<=1;
end
18'd60943: begin  
end
18'd60944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd60945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd60946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd60947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd60948: begin  
rid<=0;
end
18'd61001: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=72;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5400;
 end   
18'd61002: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=36;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=2602;
 end   
18'd61003: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=99;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=7148;
 end   
18'd61004: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=75;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=5430;
 end   
18'd61005: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=90;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=6520;
 end   
18'd61006: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=76;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=5522;
 end   
18'd61007: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=56;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=4092;
 end   
18'd61008: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd61142: begin  
rid<=1;
end
18'd61143: begin  
end
18'd61144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd61145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd61146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd61147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd61148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd61149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd61150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd61151: begin  
rid<=0;
end
18'd61201: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=42;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4239;
 end   
18'd61202: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=95;
   mapp<=15;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7365;
 end   
18'd61203: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=66;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5282;
 end   
18'd61204: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=56;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=5072;
 end   
18'd61205: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=86;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd61206: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd61207: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd61342: begin  
rid<=1;
end
18'd61343: begin  
end
18'd61344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd61345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd61346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd61347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd61348: begin  
rid<=0;
end
18'd61401: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=64;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1664;
 end   
18'd61402: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=85;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2220;
 end   
18'd61403: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=65;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1710;
 end   
18'd61404: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=8;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=238;
 end   
18'd61405: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd61542: begin  
rid<=1;
end
18'd61543: begin  
end
18'd61544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd61545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd61546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd61547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd61548: begin  
rid<=0;
end
18'd61601: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=12;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2976;
 end   
18'd61602: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=52;
   mapp<=54;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2790;
 end   
18'd61603: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=38;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=876;
 end   
18'd61604: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=6;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=1464;
 end   
18'd61605: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=25;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=2010;
 end   
18'd61606: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=30;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=3116;
 end   
18'd61607: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=49;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=5012;
 end   
18'd61608: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=79;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd61609: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd61610: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd61742: begin  
rid<=1;
end
18'd61743: begin  
end
18'd61744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd61745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd61746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd61747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd61748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd61749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd61750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd61751: begin  
rid<=0;
end
18'd61801: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=81;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14027;
 end   
18'd61802: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=70;
   mapp<=17;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=16756;
 end   
18'd61803: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=47;
   mapp<=21;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=20772;
 end   
18'd61804: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=53;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd61805: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=8;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd61806: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=8;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd61807: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=15;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd61808: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=29;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd61809: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=66;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd61810: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd61811: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd61812: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd61813: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14027;
 end   
18'd61814: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14027;
 end   
18'd61815: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14027;
 end   
18'd61816: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14027;
 end   
18'd61817: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14027;
 end   
18'd61818: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14027;
 end   
18'd61819: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14027;
 end   
18'd61820: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14027;
 end   
18'd61942: begin  
rid<=1;
end
18'd61943: begin  
end
18'd61944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd61945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd61946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd61947: begin  
rid<=0;
end
18'd62001: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=31;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2201;
 end   
18'd62002: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=41;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=1281;
 end   
18'd62003: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=59;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=1849;
 end   
18'd62004: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd62142: begin  
rid<=1;
end
18'd62143: begin  
end
18'd62144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd62145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd62146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd62147: begin  
rid<=0;
end
18'd62201: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=27;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=19102;
 end   
18'd62202: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=13;
   mapp<=88;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=19708;
 end   
18'd62203: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=23;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=15734;
 end   
18'd62204: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=71;
   mapp<=68;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=16542;
 end   
18'd62205: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=27;
   mapp<=99;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=14734;
 end   
18'd62206: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=73;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd62207: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=61;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd62208: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd62209: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd62210: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd62211: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd62212: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd62213: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19102;
 end   
18'd62214: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19102;
 end   
18'd62215: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19102;
 end   
18'd62216: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19102;
 end   
18'd62217: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19102;
 end   
18'd62218: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19102;
 end   
18'd62342: begin  
rid<=1;
end
18'd62343: begin  
end
18'd62344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd62345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd62346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd62347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd62348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd62349: begin  
rid<=0;
end
18'd62401: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=95;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1321;
 end   
18'd62402: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=13;
   mapp<=87;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8496;
 end   
18'd62403: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=17;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=2454;
 end   
18'd62404: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=63;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=6704;
 end   
18'd62405: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=53;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=5413;
 end   
18'd62406: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=26;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=3755;
 end   
18'd62407: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd62408: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd62409: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd62542: begin  
rid<=1;
end
18'd62543: begin  
end
18'd62544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd62545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd62546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd62547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd62548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd62549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd62550: begin  
rid<=0;
end
18'd62601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=93;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12152;
 end   
18'd62602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=85;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10780;
 end   
18'd62603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=65;
   mapp<=96;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=13248;
 end   
18'd62604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=33;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=8434;
 end   
18'd62605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=23;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=11734;
 end   
18'd62606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=52;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=12836;
 end   
18'd62607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=79;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=10712;
 end   
18'd62608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd62609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd62610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd62611: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd62612: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd62742: begin  
rid<=1;
end
18'd62743: begin  
end
18'd62744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd62745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd62746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd62747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd62748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd62749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd62750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd62751: begin  
rid<=0;
end
18'd62801: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=90;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=630;
 end   
18'd62802: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=71;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=6400;
 end   
18'd62803: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=87;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=7850;
 end   
18'd62804: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=99;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=8940;
 end   
18'd62805: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=19;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=1750;
 end   
18'd62806: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=96;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=8690;
 end   
18'd62807: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=15;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=1410;
 end   
18'd62808: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=52;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=4750;
 end   
18'd62809: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=92;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=8360;
 end   
18'd62810: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=53;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[9]<=4860;
 end   
18'd62811: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=57;
   pp<=100;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[10]<=5230;
 end   
18'd62812: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd62942: begin  
rid<=1;
end
18'd62943: begin  
end
18'd62944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd62945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd62946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd62947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd62948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd62949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd62950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd62951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd62952: begin  
check<=expctdoutput[8]-outcheck;
end
18'd62953: begin  
check<=expctdoutput[9]-outcheck;
end
18'd62954: begin  
check<=expctdoutput[10]-outcheck;
end
18'd62955: begin  
rid<=0;
end
18'd63001: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=9;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=774;
 end   
18'd63002: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=65;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5600;
 end   
18'd63003: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=86;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=7416;
 end   
18'd63004: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=19;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=1664;
 end   
18'd63005: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd63142: begin  
rid<=1;
end
18'd63143: begin  
end
18'd63144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd63145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd63146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd63147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd63148: begin  
rid<=0;
end
18'd63201: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=78;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13823;
 end   
18'd63202: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=74;
   mapp<=28;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=16335;
 end   
18'd63203: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=95;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd63204: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=43;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd63205: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=74;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd63206: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=16;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd63207: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd63208: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd63209: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd63210: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd63211: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd63212: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd63213: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13823;
 end   
18'd63342: begin  
rid<=1;
end
18'd63343: begin  
end
18'd63344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd63345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd63346: begin  
rid<=0;
end
18'd63401: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=22;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=19632;
 end   
18'd63402: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=83;
   mapp<=22;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=23677;
 end   
18'd63403: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=31;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd63404: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=3;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd63405: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=32;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd63406: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd63407: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=90;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd63408: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=80;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd63409: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=8;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd63410: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd63411: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd63412: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd63413: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19632;
 end   
18'd63414: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19632;
 end   
18'd63415: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19632;
 end   
18'd63416: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19632;
 end   
18'd63417: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19632;
 end   
18'd63418: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19632;
 end   
18'd63419: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19632;
 end   
18'd63542: begin  
rid<=1;
end
18'd63543: begin  
end
18'd63544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd63545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd63546: begin  
rid<=0;
end
18'd63601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=13;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16724;
 end   
18'd63602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=32;
   mapp<=18;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=18451;
 end   
18'd63603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=92;
   mapp<=57;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=19975;
 end   
18'd63604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=82;
   mapp<=61;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=19850;
 end   
18'd63605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=67;
   mapp<=20;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=21126;
 end   
18'd63606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=20;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd63607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=58;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd63608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=74;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd63609: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=87;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd63610: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=94;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd63611: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=83;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd63612: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd63613: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16724;
 end   
18'd63614: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16724;
 end   
18'd63615: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16724;
 end   
18'd63616: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16724;
 end   
18'd63617: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16724;
 end   
18'd63618: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16724;
 end   
18'd63742: begin  
rid<=1;
end
18'd63743: begin  
end
18'd63744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd63745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd63746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd63747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd63748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd63749: begin  
rid<=0;
end
18'd63801: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=25;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8550;
 end   
18'd63802: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=55;
   mapp<=46;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9708;
 end   
18'd63803: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=63;
   mapp<=90;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12264;
 end   
18'd63804: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=67;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=7990;
 end   
18'd63805: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=92;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=4464;
 end   
18'd63806: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=31;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd63807: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=19;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd63808: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd63809: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd63810: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd63942: begin  
rid<=1;
end
18'd63943: begin  
end
18'd63944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd63945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd63946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd63947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd63948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd63949: begin  
rid<=0;
end
18'd64001: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=59;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=17572;
 end   
18'd64002: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=18;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=19457;
 end   
18'd64003: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=20;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd64004: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=35;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd64005: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=14;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd64006: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=56;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd64007: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=47;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd64008: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=56;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd64009: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=34;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd64010: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=60;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd64011: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=51;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd64012: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd64013: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17572;
 end   
18'd64014: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17572;
 end   
18'd64015: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17572;
 end   
18'd64016: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17572;
 end   
18'd64017: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17572;
 end   
18'd64018: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17572;
 end   
18'd64019: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17572;
 end   
18'd64020: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17572;
 end   
18'd64021: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17572;
 end   
18'd64142: begin  
rid<=1;
end
18'd64143: begin  
end
18'd64144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd64145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd64146: begin  
rid<=0;
end
18'd64201: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=89;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=19454;
 end   
18'd64202: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=72;
   mapp<=89;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=14851;
 end   
18'd64203: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=19;
   mapp<=24;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=10959;
 end   
18'd64204: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=1;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd64205: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=2;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd64206: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=44;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd64207: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd64208: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=39;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd64209: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd64210: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd64211: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd64212: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd64213: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19454;
 end   
18'd64214: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19454;
 end   
18'd64342: begin  
rid<=1;
end
18'd64343: begin  
end
18'd64344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd64345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd64346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd64347: begin  
rid<=0;
end
18'd64401: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=14;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2512;
 end   
18'd64402: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=15;
   mapp<=86;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2642;
 end   
18'd64403: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=44;
   mapp<=16;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=3685;
 end   
18'd64404: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=27;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=2455;
 end   
18'd64405: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=69;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=5707;
 end   
18'd64406: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd64407: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd64408: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd64409: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd64410: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd64542: begin  
rid<=1;
end
18'd64543: begin  
end
18'd64544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd64545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd64546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd64547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd64548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd64549: begin  
rid<=0;
end
18'd64601: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=52;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9698;
 end   
18'd64602: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=46;
   mapp<=76;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7280;
 end   
18'd64603: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=37;
   mapp<=58;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9150;
 end   
18'd64604: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=15;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=8816;
 end   
18'd64605: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=88;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=13224;
 end   
18'd64606: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=16;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=12742;
 end   
18'd64607: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=88;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=17448;
 end   
18'd64608: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=82;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd64609: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=74;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd64610: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd64611: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd64612: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd64742: begin  
rid<=1;
end
18'd64743: begin  
end
18'd64744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd64745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd64746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd64747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd64748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd64749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd64750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd64751: begin  
rid<=0;
end
18'd64801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=42;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15362;
 end   
18'd64802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=84;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=16322;
 end   
18'd64803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=72;
   mapp<=62;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=15190;
 end   
18'd64804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=49;
   mapp<=16;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=13297;
 end   
18'd64805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=96;
   mapp<=24;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=14252;
 end   
18'd64806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=26;
   mapp<=29;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=9691;
 end   
18'd64807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=82;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd64808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=2;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd64809: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=75;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd64810: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd64811: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=65;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd64812: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd64813: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15362;
 end   
18'd64814: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15362;
 end   
18'd64815: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15362;
 end   
18'd64816: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15362;
 end   
18'd64817: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15362;
 end   
18'd64942: begin  
rid<=1;
end
18'd64943: begin  
end
18'd64944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd64945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd64946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd64947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd64948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd64949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd64950: begin  
rid<=0;
end
18'd65001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=17;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12193;
 end   
18'd65002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=93;
   mapp<=17;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=12713;
 end   
18'd65003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=73;
   mapp<=44;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=17794;
 end   
18'd65004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=60;
   mapp<=54;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=14289;
 end   
18'd65005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=75;
   mapp<=43;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=13125;
 end   
18'd65006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=24;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=15006;
 end   
18'd65007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=99;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=8277;
 end   
18'd65008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd65009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd65010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd65011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd65012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd65013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12193;
 end   
18'd65014: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12193;
 end   
18'd65015: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12193;
 end   
18'd65016: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12193;
 end   
18'd65142: begin  
rid<=1;
end
18'd65143: begin  
end
18'd65144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd65145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd65146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd65147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd65148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd65149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd65150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd65151: begin  
rid<=0;
end
18'd65201: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=93;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=269;
 end   
18'd65202: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=8;
   mapp<=22;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2120;
 end   
18'd65203: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=8;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=1524;
 end   
18'd65204: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=95;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=9073;
 end   
18'd65205: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=26;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=2618;
 end   
18'd65206: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=20;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=2638;
 end   
18'd65207: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=91;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=9227;
 end   
18'd65208: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=88;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=8486;
 end   
18'd65209: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=29;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=3353;
 end   
18'd65210: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=72;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[9]<=7402;
 end   
18'd65211: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd65212: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd65213: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=269;
 end   
18'd65342: begin  
rid<=1;
end
18'd65343: begin  
end
18'd65344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd65345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd65346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd65347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd65348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd65349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd65350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd65351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd65352: begin  
check<=expctdoutput[8]-outcheck;
end
18'd65353: begin  
check<=expctdoutput[9]-outcheck;
end
18'd65354: begin  
rid<=0;
end
18'd65401: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=37;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2812;
 end   
18'd65402: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=16;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1226;
 end   
18'd65403: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=3;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=248;
 end   
18'd65404: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=90;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=6870;
 end   
18'd65405: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=12;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=952;
 end   
18'd65406: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=89;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=6814;
 end   
18'd65407: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=53;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=4088;
 end   
18'd65408: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=79;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=6074;
 end   
18'd65409: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=99;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=7604;
 end   
18'd65410: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=22;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[9]<=1762;
 end   
18'd65411: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd65542: begin  
rid<=1;
end
18'd65543: begin  
end
18'd65544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd65545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd65546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd65547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd65548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd65549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd65550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd65551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd65552: begin  
check<=expctdoutput[8]-outcheck;
end
18'd65553: begin  
check<=expctdoutput[9]-outcheck;
end
18'd65554: begin  
rid<=0;
end
18'd65601: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=54;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3726;
 end   
18'd65602: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=29;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2011;
 end   
18'd65603: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=34;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=2366;
 end   
18'd65604: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=38;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=2652;
 end   
18'd65605: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd65742: begin  
rid<=1;
end
18'd65743: begin  
end
18'd65744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd65745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd65746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd65747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd65748: begin  
rid<=0;
end
18'd65801: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=95;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8671;
 end   
18'd65802: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=79;
   mapp<=34;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8928;
 end   
18'd65803: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=72;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=10652;
 end   
18'd65804: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=48;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=8777;
 end   
18'd65805: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=53;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=5312;
 end   
18'd65806: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=3;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=888;
 end   
18'd65807: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=7;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=2147;
 end   
18'd65808: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=18;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=4387;
 end   
18'd65809: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=33;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=6138;
 end   
18'd65810: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd65811: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd65812: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd65942: begin  
rid<=1;
end
18'd65943: begin  
end
18'd65944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd65945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd65946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd65947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd65948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd65949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd65950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd65951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd65952: begin  
check<=expctdoutput[8]-outcheck;
end
18'd65953: begin  
rid<=0;
end
18'd66001: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=7;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=413;
 end   
18'd66002: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=0;
   mapp<=61;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=437;
 end   
18'd66003: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd66142: begin  
rid<=1;
end
18'd66143: begin  
end
18'd66144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd66145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd66146: begin  
rid<=0;
end
18'd66201: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=32;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=17410;
 end   
18'd66202: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=56;
   mapp<=92;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=18730;
 end   
18'd66203: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=58;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd66204: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=49;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd66205: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=20;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd66206: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=96;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd66207: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=24;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd66208: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=20;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd66209: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=26;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd66210: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd66211: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd66212: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd66213: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17410;
 end   
18'd66214: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17410;
 end   
18'd66215: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17410;
 end   
18'd66216: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17410;
 end   
18'd66217: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17410;
 end   
18'd66218: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17410;
 end   
18'd66219: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17410;
 end   
18'd66342: begin  
rid<=1;
end
18'd66343: begin  
end
18'd66344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd66345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd66346: begin  
rid<=0;
end
18'd66401: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=4;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16021;
 end   
18'd66402: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=77;
   mapp<=74;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=15773;
 end   
18'd66403: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=53;
   mapp<=91;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=11477;
 end   
18'd66404: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=42;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd66405: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=4;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd66406: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=23;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd66407: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=52;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd66408: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=25;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd66409: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd66410: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd66411: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd66412: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd66413: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16021;
 end   
18'd66414: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16021;
 end   
18'd66542: begin  
rid<=1;
end
18'd66543: begin  
end
18'd66544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd66545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd66546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd66547: begin  
rid<=0;
end
18'd66601: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=49;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1176;
 end   
18'd66602: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=35;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=850;
 end   
18'd66603: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd66742: begin  
rid<=1;
end
18'd66743: begin  
end
18'd66744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd66745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd66746: begin  
rid<=0;
end
18'd66801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=79;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6714;
 end   
18'd66802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=2;
   mapp<=55;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11186;
 end   
18'd66803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=83;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd66804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=92;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd66805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=32;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd66806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd66807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd66808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd66809: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd66810: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd66811: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd66942: begin  
rid<=1;
end
18'd66943: begin  
end
18'd66944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd66945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd66946: begin  
rid<=0;
end
18'd67001: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=71;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=21380;
 end   
18'd67002: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=78;
   mapp<=47;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=17720;
 end   
18'd67003: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=40;
   mapp<=5;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=19779;
 end   
18'd67004: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=56;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd67005: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=48;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd67006: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=44;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd67007: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=45;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd67008: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=25;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd67009: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd67010: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd67011: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd67012: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd67013: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21380;
 end   
18'd67014: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21380;
 end   
18'd67015: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21380;
 end   
18'd67016: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21380;
 end   
18'd67017: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21380;
 end   
18'd67018: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21380;
 end   
18'd67142: begin  
rid<=1;
end
18'd67143: begin  
end
18'd67144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd67145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd67146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd67147: begin  
rid<=0;
end
18'd67201: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=79;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8704;
 end   
18'd67202: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=93;
   mapp<=80;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7725;
 end   
18'd67203: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=15;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=7157;
 end   
18'd67204: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=64;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=7504;
 end   
18'd67205: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=26;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=8790;
 end   
18'd67206: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd67207: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd67208: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd67342: begin  
rid<=1;
end
18'd67343: begin  
end
18'd67344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd67345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd67346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd67347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd67348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd67349: begin  
rid<=0;
end
18'd67401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=8;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3646;
 end   
18'd67402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=96;
   mapp<=33;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4060;
 end   
18'd67403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=38;
   mapp<=5;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9628;
 end   
18'd67404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=87;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=5242;
 end   
18'd67405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=32;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=6414;
 end   
18'd67406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=38;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=9026;
 end   
18'd67407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=65;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=7408;
 end   
18'd67408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=64;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=6072;
 end   
18'd67409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=18;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=10944;
 end   
18'd67410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd67411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd67412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd67413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=3646;
 end   
18'd67414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=3646;
 end   
18'd67542: begin  
rid<=1;
end
18'd67543: begin  
end
18'd67544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd67545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd67546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd67547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd67548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd67549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd67550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd67551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd67552: begin  
check<=expctdoutput[8]-outcheck;
end
18'd67553: begin  
rid<=0;
end
18'd67601: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=43;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1935;
 end   
18'd67602: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=59;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=2547;
 end   
18'd67603: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=69;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=2987;
 end   
18'd67604: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=44;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=1922;
 end   
18'd67605: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=62;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=2706;
 end   
18'd67606: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=69;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=3017;
 end   
18'd67607: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=49;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=2167;
 end   
18'd67608: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=18;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=844;
 end   
18'd67609: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=67;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=2961;
 end   
18'd67610: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=58;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[9]<=2584;
 end   
18'd67611: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd67742: begin  
rid<=1;
end
18'd67743: begin  
end
18'd67744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd67745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd67746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd67747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd67748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd67749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd67750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd67751: begin  
check<=expctdoutput[7]-outcheck;
end
18'd67752: begin  
check<=expctdoutput[8]-outcheck;
end
18'd67753: begin  
check<=expctdoutput[9]-outcheck;
end
18'd67754: begin  
rid<=0;
end
18'd67801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=68;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9872;
 end   
18'd67802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=23;
   mapp<=86;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8936;
 end   
18'd67803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=47;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd67804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=96;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd67805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=66;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd67806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=30;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd67807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=65;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd67808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd67809: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd67810: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd67811: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd67812: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd67813: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9872;
 end   
18'd67942: begin  
rid<=1;
end
18'd67943: begin  
end
18'd67944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd67945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd67946: begin  
rid<=0;
end
18'd68001: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=24;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2452;
 end   
18'd68002: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=28;
   mapp<=73;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4170;
 end   
18'd68003: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=86;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=3988;
 end   
18'd68004: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=68;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=4378;
 end   
18'd68005: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=97;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=4580;
 end   
18'd68006: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd68007: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd68008: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd68142: begin  
rid<=1;
end
18'd68143: begin  
end
18'd68144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd68145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd68146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd68147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd68148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd68149: begin  
rid<=0;
end
18'd68201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=52;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9047;
 end   
18'd68202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=69;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd68203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=62;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd68204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=70;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd68205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd68206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd68207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd68208: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd68342: begin  
rid<=1;
end
18'd68343: begin  
end
18'd68344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd68345: begin  
rid<=0;
end
18'd68401: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=67;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=18832;
 end   
18'd68402: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=54;
   mapp<=11;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=16645;
 end   
18'd68403: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=87;
   mapp<=64;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=22862;
 end   
18'd68404: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=17;
   mapp<=50;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=14418;
 end   
18'd68405: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=65;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd68406: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=42;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd68407: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd68408: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=73;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd68409: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=15;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd68410: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd68411: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd68412: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd68413: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18832;
 end   
18'd68414: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18832;
 end   
18'd68415: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18832;
 end   
18'd68542: begin  
rid<=1;
end
18'd68543: begin  
end
18'd68544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd68545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd68546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd68547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd68548: begin  
rid<=0;
end
18'd68601: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=30;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6701;
 end   
18'd68602: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=9;
   mapp<=69;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5368;
 end   
18'd68603: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=40;
   mapp<=86;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6623;
 end   
18'd68604: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=21;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd68605: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=19;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd68606: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd68607: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd68608: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd68742: begin  
rid<=1;
end
18'd68743: begin  
end
18'd68744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd68745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd68746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd68747: begin  
rid<=0;
end
18'd68801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=99;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2376;
 end   
18'd68802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=36;
   mapp<=11;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3043;
 end   
18'd68803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=54;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=8714;
 end   
18'd68804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=93;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=12261;
 end   
18'd68805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=84;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=10408;
 end   
18'd68806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd68807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd68808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd68942: begin  
rid<=1;
end
18'd68943: begin  
end
18'd68944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd68945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd68946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd68947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd68948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd68949: begin  
rid<=0;
end
18'd69001: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=17;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=20369;
 end   
18'd69002: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=13;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=20573;
 end   
18'd69003: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=53;
   mapp<=65;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=29554;
 end   
18'd69004: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=17;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd69005: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=77;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd69006: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=60;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd69007: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=5;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd69008: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=53;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd69009: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=91;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd69010: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd69011: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=76;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd69012: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd69013: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20369;
 end   
18'd69014: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20369;
 end   
18'd69015: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20369;
 end   
18'd69016: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20369;
 end   
18'd69017: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20369;
 end   
18'd69018: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20369;
 end   
18'd69019: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20369;
 end   
18'd69020: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20369;
 end   
18'd69142: begin  
rid<=1;
end
18'd69143: begin  
end
18'd69144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd69145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd69146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd69147: begin  
rid<=0;
end
18'd69201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=45;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6665;
 end   
18'd69202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=52;
   mapp<=16;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9253;
 end   
18'd69203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=47;
   mapp<=50;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9096;
 end   
18'd69204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=21;
   mapp<=93;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=9407;
 end   
18'd69205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=61;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=11906;
 end   
18'd69206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=44;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=13695;
 end   
18'd69207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=59;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd69208: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=66;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd69209: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=85;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd69210: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd69211: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd69212: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd69213: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6665;
 end   
18'd69342: begin  
rid<=1;
end
18'd69343: begin  
end
18'd69344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd69345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd69346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd69347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd69348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd69349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd69350: begin  
rid<=0;
end
18'd69401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=98;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6942;
 end   
18'd69402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=92;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11642;
 end   
18'd69403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=54;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=9912;
 end   
18'd69404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=50;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=7874;
 end   
18'd69405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=32;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=12284;
 end   
18'd69406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=99;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=11592;
 end   
18'd69407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=20;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=5240;
 end   
18'd69408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd69409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd69410: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd69542: begin  
rid<=1;
end
18'd69543: begin  
end
18'd69544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd69545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd69546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd69547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd69548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd69549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd69550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd69551: begin  
rid<=0;
end
18'd69601: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=16;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=464;
 end   
18'd69602: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=59;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1721;
 end   
18'd69603: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=58;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1702;
 end   
18'd69604: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd69742: begin  
rid<=1;
end
18'd69743: begin  
end
18'd69744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd69745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd69746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd69747: begin  
rid<=0;
end
18'd69801: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=95;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12129;
 end   
18'd69802: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=86;
   mapp<=57;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13842;
 end   
18'd69803: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=3;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=17062;
 end   
18'd69804: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=52;
   mapp<=71;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=14631;
 end   
18'd69805: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=42;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=11453;
 end   
18'd69806: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd69807: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd69808: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd69809: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd69810: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd69811: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd69812: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd69942: begin  
rid<=1;
end
18'd69943: begin  
end
18'd69944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd69945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd69946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd69947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd69948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd69949: begin  
rid<=0;
end
18'd70001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=41;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4549;
 end   
18'd70002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=38;
   mapp<=28;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4122;
 end   
18'd70003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=78;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=5498;
 end   
18'd70004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=60;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=2528;
 end   
18'd70005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=1;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=1943;
 end   
18'd70006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=49;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=4491;
 end   
18'd70007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=64;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=5914;
 end   
18'd70008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=85;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=4543;
 end   
18'd70009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=26;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=3312;
 end   
18'd70010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=57;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[9]<=3833;
 end   
18'd70011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd70012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd70013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=4549;
 end   
18'd70142: begin  
rid<=1;
end
18'd70143: begin  
end
18'd70144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd70145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd70146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd70147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd70148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd70149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd70150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd70151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd70152: begin  
check<=expctdoutput[8]-outcheck;
end
18'd70153: begin  
check<=expctdoutput[9]-outcheck;
end
18'd70154: begin  
rid<=0;
end
18'd70201: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=23;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12074;
 end   
18'd70202: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=99;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11144;
 end   
18'd70203: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=31;
   mapp<=68;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9896;
 end   
18'd70204: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=73;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=5453;
 end   
18'd70205: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=35;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=4712;
 end   
18'd70206: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=9;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=12272;
 end   
18'd70207: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=96;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=12178;
 end   
18'd70208: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=81;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=9181;
 end   
18'd70209: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=61;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=7948;
 end   
18'd70210: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd70211: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd70212: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd70213: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12074;
 end   
18'd70214: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12074;
 end   
18'd70342: begin  
rid<=1;
end
18'd70343: begin  
end
18'd70344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd70345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd70346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd70347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd70348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd70349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd70350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd70351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd70352: begin  
check<=expctdoutput[8]-outcheck;
end
18'd70353: begin  
rid<=0;
end
18'd70401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=40;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5691;
 end   
18'd70402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=69;
   mapp<=50;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9230;
 end   
18'd70403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=23;
   mapp<=87;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=10387;
 end   
18'd70404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=88;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=11129;
 end   
18'd70405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=67;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=4592;
 end   
18'd70406: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=83;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=5594;
 end   
18'd70407: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=3482;
 end   
18'd70408: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=58;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=4024;
 end   
18'd70409: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=6;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=7497;
 end   
18'd70410: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd70411: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=63;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd70412: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd70413: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5691;
 end   
18'd70414: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5691;
 end   
18'd70542: begin  
rid<=1;
end
18'd70543: begin  
end
18'd70544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd70545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd70546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd70547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd70548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd70549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd70550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd70551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd70552: begin  
check<=expctdoutput[8]-outcheck;
end
18'd70553: begin  
rid<=0;
end
18'd70601: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=88;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=26006;
 end   
18'd70602: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=19;
   mapp<=85;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=32472;
 end   
18'd70603: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=46;
   mapp<=23;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=27795;
 end   
18'd70604: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=90;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd70605: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=75;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd70606: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=69;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd70607: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=19;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd70608: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=41;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd70609: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd70610: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd70611: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd70612: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd70613: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26006;
 end   
18'd70614: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26006;
 end   
18'd70615: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26006;
 end   
18'd70616: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26006;
 end   
18'd70617: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26006;
 end   
18'd70618: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26006;
 end   
18'd70742: begin  
rid<=1;
end
18'd70743: begin  
end
18'd70744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd70745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd70746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd70747: begin  
rid<=0;
end
18'd70801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=18386;
 end   
18'd70802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=32;
   mapp<=58;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=23451;
 end   
18'd70803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=75;
   mapp<=58;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=25060;
 end   
18'd70804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=36;
   mapp<=94;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=26438;
 end   
18'd70805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=38;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd70806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=58;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd70807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=80;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd70808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=85;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd70809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=13;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd70810: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=84;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd70811: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd70812: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd70813: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18386;
 end   
18'd70814: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18386;
 end   
18'd70815: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18386;
 end   
18'd70816: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18386;
 end   
18'd70817: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18386;
 end   
18'd70942: begin  
rid<=1;
end
18'd70943: begin  
end
18'd70944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd70945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd70946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd70947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd70948: begin  
rid<=0;
end
18'd71001: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=48;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14272;
 end   
18'd71002: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=77;
   mapp<=26;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13047;
 end   
18'd71003: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=99;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=16621;
 end   
18'd71004: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=35;
   mapp<=36;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=16640;
 end   
18'd71005: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd71006: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd71007: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd71008: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd71009: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd71010: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd71011: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd71142: begin  
rid<=1;
end
18'd71143: begin  
end
18'd71144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd71145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd71146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd71147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd71148: begin  
rid<=0;
end
18'd71201: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=67;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=21782;
 end   
18'd71202: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=31;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=20038;
 end   
18'd71203: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=28;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd71204: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=16;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd71205: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=34;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd71206: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=99;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd71207: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=57;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd71208: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=40;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd71209: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=81;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd71210: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=23;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd71211: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=41;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd71212: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd71213: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21782;
 end   
18'd71214: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21782;
 end   
18'd71215: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21782;
 end   
18'd71216: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21782;
 end   
18'd71217: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21782;
 end   
18'd71218: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21782;
 end   
18'd71219: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21782;
 end   
18'd71220: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21782;
 end   
18'd71221: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21782;
 end   
18'd71342: begin  
rid<=1;
end
18'd71343: begin  
end
18'd71344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd71345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd71346: begin  
rid<=0;
end
18'd71401: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=63;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8961;
 end   
18'd71402: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=45;
   mapp<=99;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6790;
 end   
18'd71403: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=26;
   mapp<=75;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=11150;
 end   
18'd71404: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=1;
   mapp<=99;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=17481;
 end   
18'd71405: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=24;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=19333;
 end   
18'd71406: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=83;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=17099;
 end   
18'd71407: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd71408: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=35;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd71409: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=24;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd71410: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd71411: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd71412: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd71413: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8961;
 end   
18'd71542: begin  
rid<=1;
end
18'd71543: begin  
end
18'd71544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd71545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd71546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd71547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd71548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd71549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd71550: begin  
rid<=0;
end
18'd71601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=68;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11301;
 end   
18'd71602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=70;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10800;
 end   
18'd71603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=43;
   mapp<=17;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9852;
 end   
18'd71604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=92;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=10958;
 end   
18'd71605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=52;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=8395;
 end   
18'd71606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=24;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=8512;
 end   
18'd71607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=73;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=10189;
 end   
18'd71608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd71609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd71610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd71611: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd71612: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd71742: begin  
rid<=1;
end
18'd71743: begin  
end
18'd71744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd71745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd71746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd71747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd71748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd71749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd71750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd71751: begin  
rid<=0;
end
18'd71801: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=28;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=19700;
 end   
18'd71802: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=90;
   mapp<=14;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=19664;
 end   
18'd71803: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=99;
   mapp<=80;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=15702;
 end   
18'd71804: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=80;
   mapp<=58;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=10660;
 end   
18'd71805: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=70;
   mapp<=58;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=10186;
 end   
18'd71806: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=24;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=9081;
 end   
18'd71807: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd71808: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd71809: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd71810: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd71811: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd71812: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd71813: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19700;
 end   
18'd71814: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19700;
 end   
18'd71815: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19700;
 end   
18'd71942: begin  
rid<=1;
end
18'd71943: begin  
end
18'd71944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd71945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd71946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd71947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd71948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd71949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd71950: begin  
rid<=0;
end
18'd72001: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=36;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11124;
 end   
18'd72002: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=66;
   mapp<=64;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=14992;
 end   
18'd72003: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=92;
   mapp<=75;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=15808;
 end   
18'd72004: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=84;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=9478;
 end   
18'd72005: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=82;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=4270;
 end   
18'd72006: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=11;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=7098;
 end   
18'd72007: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=6;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=8812;
 end   
18'd72008: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=68;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=7814;
 end   
18'd72009: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd72010: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd72011: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd72012: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd72013: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11124;
 end   
18'd72142: begin  
rid<=1;
end
18'd72143: begin  
end
18'd72144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd72145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd72146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd72147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd72148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd72149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd72150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd72151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd72152: begin  
rid<=0;
end
18'd72201: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=10;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14981;
 end   
18'd72202: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=57;
   mapp<=12;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=17030;
 end   
18'd72203: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=66;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd72204: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=50;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd72205: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=70;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd72206: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=45;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd72207: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=25;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd72208: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd72209: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd72210: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd72211: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd72212: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd72213: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14981;
 end   
18'd72214: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14981;
 end   
18'd72215: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14981;
 end   
18'd72342: begin  
rid<=1;
end
18'd72343: begin  
end
18'd72344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd72345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd72346: begin  
rid<=0;
end
18'd72401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=1;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=74;
 end   
18'd72402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=43;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=53;
 end   
18'd72403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=29;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=49;
 end   
18'd72404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=36;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=66;
 end   
18'd72405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=63;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=103;
 end   
18'd72406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=16;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=66;
 end   
18'd72407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=58;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=118;
 end   
18'd72408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=34;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=104;
 end   
18'd72409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd72542: begin  
rid<=1;
end
18'd72543: begin  
end
18'd72544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd72545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd72546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd72547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd72548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd72549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd72550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd72551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd72552: begin  
rid<=0;
end
18'd72601: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=24;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14185;
 end   
18'd72602: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=74;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11558;
 end   
18'd72603: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=75;
   mapp<=82;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12083;
 end   
18'd72604: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=37;
   mapp<=39;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=12393;
 end   
18'd72605: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=76;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd72606: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd72607: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=24;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd72608: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=64;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd72609: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd72610: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd72611: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd72612: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd72613: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14185;
 end   
18'd72742: begin  
rid<=1;
end
18'd72743: begin  
end
18'd72744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd72745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd72746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd72747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd72748: begin  
rid<=0;
end
18'd72801: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=29;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=725;
 end   
18'd72802: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd72942: begin  
rid<=1;
end
18'd72943: begin  
end
18'd72944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd72945: begin  
rid<=0;
end
18'd73001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=90;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8460;
 end   
18'd73002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=44;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=3970;
 end   
18'd73003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=6;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=560;
 end   
18'd73004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=75;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=6780;
 end   
18'd73005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=71;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=6430;
 end   
18'd73006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd73142: begin  
rid<=1;
end
18'd73143: begin  
end
18'd73144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd73145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd73146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd73147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd73148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd73149: begin  
rid<=0;
end
18'd73201: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=56;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8180;
 end   
18'd73202: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=20;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6714;
 end   
18'd73203: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=32;
   mapp<=58;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=4848;
 end   
18'd73204: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=7;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=3690;
 end   
18'd73205: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=45;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=5256;
 end   
18'd73206: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd73207: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd73208: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd73209: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd73210: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd73342: begin  
rid<=1;
end
18'd73343: begin  
end
18'd73344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd73345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd73346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd73347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd73348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd73349: begin  
rid<=0;
end
18'd73401: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=94;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=23565;
 end   
18'd73402: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=90;
   mapp<=53;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=24759;
 end   
18'd73403: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=48;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd73404: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=54;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd73405: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=17;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd73406: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=92;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd73407: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=30;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd73408: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=18;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd73409: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=48;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd73410: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd73411: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd73412: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd73413: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23565;
 end   
18'd73414: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23565;
 end   
18'd73415: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23565;
 end   
18'd73416: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23565;
 end   
18'd73417: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23565;
 end   
18'd73418: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23565;
 end   
18'd73419: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23565;
 end   
18'd73542: begin  
rid<=1;
end
18'd73543: begin  
end
18'd73544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd73545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd73546: begin  
rid<=0;
end
18'd73601: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=35;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2870;
 end   
18'd73602: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=43;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=1515;
 end   
18'd73603: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=39;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=1385;
 end   
18'd73604: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=1;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=65;
 end   
18'd73605: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=93;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=3295;
 end   
18'd73606: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=27;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=995;
 end   
18'd73607: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=69;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=2475;
 end   
18'd73608: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=93;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=3325;
 end   
18'd73609: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=33;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=1235;
 end   
18'd73610: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=31;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[9]<=1175;
 end   
18'd73611: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=92;
   pp<=100;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[10]<=3320;
 end   
18'd73612: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd73742: begin  
rid<=1;
end
18'd73743: begin  
end
18'd73744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd73745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd73746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd73747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd73748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd73749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd73750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd73751: begin  
check<=expctdoutput[7]-outcheck;
end
18'd73752: begin  
check<=expctdoutput[8]-outcheck;
end
18'd73753: begin  
check<=expctdoutput[9]-outcheck;
end
18'd73754: begin  
check<=expctdoutput[10]-outcheck;
end
18'd73755: begin  
rid<=0;
end
18'd73801: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=21;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2992;
 end   
18'd73802: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=82;
   mapp<=16;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5348;
 end   
18'd73803: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=61;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=2695;
 end   
18'd73804: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=17;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=961;
 end   
18'd73805: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=7;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=1827;
 end   
18'd73806: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=20;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=4160;
 end   
18'd73807: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=45;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=6417;
 end   
18'd73808: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd73809: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd73810: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd73942: begin  
rid<=1;
end
18'd73943: begin  
end
18'd73944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd73945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd73946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd73947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd73948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd73949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd73950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd73951: begin  
rid<=0;
end
18'd74001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=81;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12061;
 end   
18'd74002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=67;
   mapp<=70;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6685;
 end   
18'd74003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=15;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=7600;
 end   
18'd74004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=95;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=10606;
 end   
18'd74005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=43;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=7744;
 end   
18'd74006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=63;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=9910;
 end   
18'd74007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=71;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=11975;
 end   
18'd74008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=92;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=9867;
 end   
18'd74009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=35;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=4054;
 end   
18'd74010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=17;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[9]<=2271;
 end   
18'd74011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd74012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd74013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12061;
 end   
18'd74142: begin  
rid<=1;
end
18'd74143: begin  
end
18'd74144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd74145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd74146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd74147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd74148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd74149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd74150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd74151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd74152: begin  
check<=expctdoutput[8]-outcheck;
end
18'd74153: begin  
check<=expctdoutput[9]-outcheck;
end
18'd74154: begin  
rid<=0;
end
18'd74201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=29;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1310;
 end   
18'd74202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=24;
   mapp<=28;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1542;
 end   
18'd74203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd74204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd74205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd74342: begin  
rid<=1;
end
18'd74343: begin  
end
18'd74344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd74345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd74346: begin  
rid<=0;
end
18'd74401: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=94;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4794;
 end   
18'd74402: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=41;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2101;
 end   
18'd74403: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=64;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=3284;
 end   
18'd74404: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=83;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=4263;
 end   
18'd74405: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=20;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=1060;
 end   
18'd74406: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=44;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=2294;
 end   
18'd74407: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=88;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=4548;
 end   
18'd74408: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=77;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=3997;
 end   
18'd74409: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd74542: begin  
rid<=1;
end
18'd74543: begin  
end
18'd74544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd74545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd74546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd74547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd74548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd74549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd74550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd74551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd74552: begin  
rid<=0;
end
18'd74601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=95;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=21846;
 end   
18'd74602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=1;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=16087;
 end   
18'd74603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=5;
   mapp<=53;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=13738;
 end   
18'd74604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=58;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd74605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=23;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd74606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=87;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd74607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=41;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd74608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=26;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd74609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=30;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd74610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=9;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd74611: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=20;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd74612: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd74613: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21846;
 end   
18'd74614: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21846;
 end   
18'd74615: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21846;
 end   
18'd74616: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21846;
 end   
18'd74617: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21846;
 end   
18'd74618: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21846;
 end   
18'd74619: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21846;
 end   
18'd74620: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21846;
 end   
18'd74742: begin  
rid<=1;
end
18'd74743: begin  
end
18'd74744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd74745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd74746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd74747: begin  
rid<=0;
end
18'd74801: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=74;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2294;
 end   
18'd74802: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=2;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=72;
 end   
18'd74803: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=20;
 end   
18'd74804: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=71;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=2231;
 end   
18'd74805: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd74942: begin  
rid<=1;
end
18'd74943: begin  
end
18'd74944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd74945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd74946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd74947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd74948: begin  
rid<=0;
end
18'd75001: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=88;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13450;
 end   
18'd75002: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=55;
   mapp<=94;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=18231;
 end   
18'd75003: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=60;
   mapp<=22;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=13475;
 end   
18'd75004: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=45;
   mapp<=36;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=16074;
 end   
18'd75005: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=23;
   mapp<=90;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=17607;
 end   
18'd75006: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=42;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd75007: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd75008: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd75009: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd75010: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd75011: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd75012: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd75013: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13450;
 end   
18'd75014: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13450;
 end   
18'd75015: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13450;
 end   
18'd75016: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13450;
 end   
18'd75142: begin  
rid<=1;
end
18'd75143: begin  
end
18'd75144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd75145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd75146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd75147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd75148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd75149: begin  
rid<=0;
end
18'd75201: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=79;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=24360;
 end   
18'd75202: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=7;
   mapp<=47;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=23872;
 end   
18'd75203: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=13;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd75204: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=60;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd75205: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=47;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd75206: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=46;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd75207: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=71;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd75208: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd75209: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd75210: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd75211: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd75212: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd75213: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24360;
 end   
18'd75214: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24360;
 end   
18'd75215: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24360;
 end   
18'd75342: begin  
rid<=1;
end
18'd75343: begin  
end
18'd75344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd75345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd75346: begin  
rid<=0;
end
18'd75401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=51;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7866;
 end   
18'd75402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=90;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7765;
 end   
18'd75403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=39;
   mapp<=36;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8537;
 end   
18'd75404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=53;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=10575;
 end   
18'd75405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=49;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=11356;
 end   
18'd75406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=88;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=7583;
 end   
18'd75407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd75408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd75409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd75410: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd75411: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd75542: begin  
rid<=1;
end
18'd75543: begin  
end
18'd75544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd75545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd75546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd75547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd75548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd75549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd75550: begin  
rid<=0;
end
18'd75601: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=3;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12425;
 end   
18'd75602: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=81;
   mapp<=24;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=15913;
 end   
18'd75603: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=77;
   mapp<=78;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=16689;
 end   
18'd75604: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=50;
   mapp<=85;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=18382;
 end   
18'd75605: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=48;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=14012;
 end   
18'd75606: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd75607: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=94;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd75608: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd75609: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd75610: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd75611: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd75612: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd75742: begin  
rid<=1;
end
18'd75743: begin  
end
18'd75744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd75745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd75746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd75747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd75748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd75749: begin  
rid<=0;
end
18'd75801: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=52;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4418;
 end   
18'd75802: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=62;
   mapp<=15;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7505;
 end   
18'd75803: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=21;
   mapp<=72;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=3839;
 end   
18'd75804: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=67;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd75805: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=28;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd75806: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd75807: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd75808: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd75942: begin  
rid<=1;
end
18'd75943: begin  
end
18'd75944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd75945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd75946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd75947: begin  
rid<=0;
end
18'd76001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=35;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15586;
 end   
18'd76002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=40;
   mapp<=82;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=18358;
 end   
18'd76003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=66;
   mapp<=89;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=16052;
 end   
18'd76004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=32;
   mapp<=86;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=12263;
 end   
18'd76005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=85;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd76006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=22;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd76007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=3;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd76008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=61;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd76009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd76010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd76011: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd76012: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd76013: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15586;
 end   
18'd76142: begin  
rid<=1;
end
18'd76143: begin  
end
18'd76144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd76145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd76146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd76147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd76148: begin  
rid<=0;
end
18'd76201: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=65;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9610;
 end   
18'd76202: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=45;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd76203: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=20;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd76204: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=10;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd76205: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=28;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd76206: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=70;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd76207: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd76208: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd76209: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd76210: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd76211: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd76212: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd76342: begin  
rid<=1;
end
18'd76343: begin  
end
18'd76344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd76345: begin  
rid<=0;
end
18'd76401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=61;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=26180;
 end   
18'd76402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=95;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd76403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=51;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd76404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=66;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd76405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=83;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd76406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=10;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd76407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=58;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd76408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=72;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd76409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=95;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd76410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=6;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd76411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=14;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd76412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd76413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26180;
 end   
18'd76414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26180;
 end   
18'd76415: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26180;
 end   
18'd76416: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26180;
 end   
18'd76417: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26180;
 end   
18'd76418: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26180;
 end   
18'd76419: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26180;
 end   
18'd76420: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26180;
 end   
18'd76421: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26180;
 end   
18'd76422: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26180;
 end   
18'd76542: begin  
rid<=1;
end
18'd76543: begin  
end
18'd76544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd76545: begin  
rid<=0;
end
18'd76601: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=87;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=435;
 end   
18'd76602: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=12;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=1054;
 end   
18'd76603: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=21;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=1847;
 end   
18'd76604: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=41;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=3597;
 end   
18'd76605: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=75;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=6565;
 end   
18'd76606: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=90;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=7880;
 end   
18'd76607: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=25;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=2235;
 end   
18'd76608: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=11;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=1027;
 end   
18'd76609: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=67;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=5909;
 end   
18'd76610: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=82;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[9]<=7224;
 end   
18'd76611: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=83;
   pp<=100;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[10]<=7321;
 end   
18'd76612: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd76742: begin  
rid<=1;
end
18'd76743: begin  
end
18'd76744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd76745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd76746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd76747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd76748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd76749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd76750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd76751: begin  
check<=expctdoutput[7]-outcheck;
end
18'd76752: begin  
check<=expctdoutput[8]-outcheck;
end
18'd76753: begin  
check<=expctdoutput[9]-outcheck;
end
18'd76754: begin  
check<=expctdoutput[10]-outcheck;
end
18'd76755: begin  
rid<=0;
end
18'd76801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=5;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=395;
 end   
18'd76802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=350;
 end   
18'd76803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=74;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=390;
 end   
18'd76804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=84;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=450;
 end   
18'd76805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=29;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=185;
 end   
18'd76806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=35;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=225;
 end   
18'd76807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=60;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=360;
 end   
18'd76808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd76942: begin  
rid<=1;
end
18'd76943: begin  
end
18'd76944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd76945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd76946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd76947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd76948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd76949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd76950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd76951: begin  
rid<=0;
end
18'd77001: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=23;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=552;
 end   
18'd77002: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=50;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=1160;
 end   
18'd77003: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=16;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=388;
 end   
18'd77004: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=60;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=1410;
 end   
18'd77005: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=1;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=63;
 end   
18'd77006: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=59;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=1407;
 end   
18'd77007: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=9;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=267;
 end   
18'd77008: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd77142: begin  
rid<=1;
end
18'd77143: begin  
end
18'd77144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd77145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd77146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd77147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd77148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd77149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd77150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd77151: begin  
rid<=0;
end
18'd77201: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=40;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3688;
 end   
18'd77202: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=48;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4290;
 end   
18'd77203: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=55;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1787;
 end   
18'd77204: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=7;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=2949;
 end   
18'd77205: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=49;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=6361;
 end   
18'd77206: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=91;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=5685;
 end   
18'd77207: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=60;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=6152;
 end   
18'd77208: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=82;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd77209: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd77210: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd77342: begin  
rid<=1;
end
18'd77343: begin  
end
18'd77344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd77345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd77346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd77347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd77348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd77349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd77350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd77351: begin  
rid<=0;
end
18'd77401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=7;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2490;
 end   
18'd77402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=25;
   mapp<=79;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1207;
 end   
18'd77403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=1;
   mapp<=25;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=679;
 end   
18'd77404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=19;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=389;
 end   
18'd77405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=9;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=159;
 end   
18'd77406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=1;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=856;
 end   
18'd77407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd77408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd77409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd77410: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd77411: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd77542: begin  
rid<=1;
end
18'd77543: begin  
end
18'd77544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd77545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd77546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd77547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd77548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd77549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd77550: begin  
rid<=0;
end
18'd77601: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=64;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5632;
 end   
18'd77602: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=63;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5554;
 end   
18'd77603: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=24;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=2132;
 end   
18'd77604: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=34;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=3022;
 end   
18'd77605: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=70;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=6200;
 end   
18'd77606: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=51;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=4538;
 end   
18'd77607: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=97;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=8596;
 end   
18'd77608: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=24;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=2182;
 end   
18'd77609: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=11;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=1048;
 end   
18'd77610: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=67;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[9]<=5986;
 end   
18'd77611: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd77742: begin  
rid<=1;
end
18'd77743: begin  
end
18'd77744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd77745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd77746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd77747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd77748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd77749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd77750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd77751: begin  
check<=expctdoutput[7]-outcheck;
end
18'd77752: begin  
check<=expctdoutput[8]-outcheck;
end
18'd77753: begin  
check<=expctdoutput[9]-outcheck;
end
18'd77754: begin  
rid<=0;
end
18'd77801: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=27;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11735;
 end   
18'd77802: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=60;
   mapp<=55;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=12536;
 end   
18'd77803: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=39;
   mapp<=28;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12231;
 end   
18'd77804: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=66;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd77805: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=37;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd77806: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=48;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd77807: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=48;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd77808: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd77809: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd77810: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd77811: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd77812: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd77942: begin  
rid<=1;
end
18'd77943: begin  
end
18'd77944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd77945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd77946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd77947: begin  
rid<=0;
end
18'd78001: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=62;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=18342;
 end   
18'd78002: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=54;
   mapp<=21;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=17421;
 end   
18'd78003: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=76;
   mapp<=33;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=17361;
 end   
18'd78004: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=54;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd78005: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=58;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd78006: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=21;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd78007: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=84;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd78008: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd78009: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=66;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd78010: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd78011: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd78012: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd78013: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18342;
 end   
18'd78014: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18342;
 end   
18'd78015: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18342;
 end   
18'd78016: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18342;
 end   
18'd78142: begin  
rid<=1;
end
18'd78143: begin  
end
18'd78144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd78145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd78146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd78147: begin  
rid<=0;
end
18'd78201: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=37;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3801;
 end   
18'd78202: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=29;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd78203: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd78204: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd78342: begin  
rid<=1;
end
18'd78343: begin  
end
18'd78344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd78345: begin  
rid<=0;
end
18'd78401: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=66;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=28295;
 end   
18'd78402: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=72;
   mapp<=1;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=29034;
 end   
18'd78403: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=93;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd78404: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=58;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd78405: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=79;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd78406: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=83;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd78407: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=87;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd78408: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=23;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd78409: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=97;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd78410: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=96;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd78411: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd78412: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd78413: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28295;
 end   
18'd78414: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28295;
 end   
18'd78415: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28295;
 end   
18'd78416: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28295;
 end   
18'd78417: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28295;
 end   
18'd78418: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28295;
 end   
18'd78419: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28295;
 end   
18'd78542: begin  
rid<=1;
end
18'd78543: begin  
end
18'd78544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd78545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd78546: begin  
rid<=0;
end
18'd78601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=24;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2103;
 end   
18'd78602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=33;
   mapp<=20;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4693;
 end   
18'd78603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=57;
   mapp<=3;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=3608;
 end   
18'd78604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=72;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=4242;
 end   
18'd78605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=20;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=4597;
 end   
18'd78606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd78607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd78608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd78609: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd78610: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd78742: begin  
rid<=1;
end
18'd78743: begin  
end
18'd78744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd78745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd78746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd78747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd78748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd78749: begin  
rid<=0;
end
18'd78801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=66;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11310;
 end   
18'd78802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=90;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11766;
 end   
18'd78803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=68;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=7202;
 end   
18'd78804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=26;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=3986;
 end   
18'd78805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=28;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd78806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd78807: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd78942: begin  
rid<=1;
end
18'd78943: begin  
end
18'd78944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd78945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd78946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd78947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd78948: begin  
rid<=0;
end
18'd79001: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=27;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13244;
 end   
18'd79002: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=82;
   mapp<=49;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=14266;
 end   
18'd79003: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=93;
   mapp<=33;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12991;
 end   
18'd79004: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=87;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd79005: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=63;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd79006: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=61;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd79007: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=65;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd79008: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=99;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd79009: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=51;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd79010: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=18;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd79011: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd79012: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd79013: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13244;
 end   
18'd79014: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13244;
 end   
18'd79015: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13244;
 end   
18'd79016: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13244;
 end   
18'd79017: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13244;
 end   
18'd79018: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13244;
 end   
18'd79142: begin  
rid<=1;
end
18'd79143: begin  
end
18'd79144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd79145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd79146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd79147: begin  
rid<=0;
end
18'd79201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=64;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7872;
 end   
18'd79202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=57;
   mapp<=58;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6871;
 end   
18'd79203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=72;
   mapp<=38;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6658;
 end   
18'd79204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=21;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd79205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=22;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd79206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=56;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd79207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd79208: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd79209: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd79210: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd79342: begin  
rid<=1;
end
18'd79343: begin  
end
18'd79344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd79345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd79346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd79347: begin  
rid<=0;
end
18'd79401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=81;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=26859;
 end   
18'd79402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=51;
   mapp<=43;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=21058;
 end   
18'd79403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=60;
   mapp<=34;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=24986;
 end   
18'd79404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=98;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd79405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=71;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd79406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=42;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd79407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=94;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd79408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=84;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd79409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=35;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd79410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd79411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd79412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd79413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26859;
 end   
18'd79414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26859;
 end   
18'd79415: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26859;
 end   
18'd79416: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26859;
 end   
18'd79417: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26859;
 end   
18'd79418: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26859;
 end   
18'd79419: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26859;
 end   
18'd79420: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26859;
 end   
18'd79542: begin  
rid<=1;
end
18'd79543: begin  
end
18'd79544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd79545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd79546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd79547: begin  
rid<=0;
end
18'd79601: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=23;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1265;
 end   
18'd79602: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=50;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2760;
 end   
18'd79603: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=88;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=4860;
 end   
18'd79604: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=39;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=2175;
 end   
18'd79605: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=10;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=590;
 end   
18'd79606: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=17;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=985;
 end   
18'd79607: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=32;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=1820;
 end   
18'd79608: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=48;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=2710;
 end   
18'd79609: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=10;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=630;
 end   
18'd79610: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=95;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[9]<=5315;
 end   
18'd79611: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=19;
   mapp<=0;
   pp<=100;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[10]<=1145;
 end   
18'd79612: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd79742: begin  
rid<=1;
end
18'd79743: begin  
end
18'd79744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd79745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd79746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd79747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd79748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd79749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd79750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd79751: begin  
check<=expctdoutput[7]-outcheck;
end
18'd79752: begin  
check<=expctdoutput[8]-outcheck;
end
18'd79753: begin  
check<=expctdoutput[9]-outcheck;
end
18'd79754: begin  
check<=expctdoutput[10]-outcheck;
end
18'd79755: begin  
rid<=0;
end
18'd79801: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=34;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16436;
 end   
18'd79802: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=84;
   mapp<=51;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=17095;
 end   
18'd79803: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=77;
   mapp<=95;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=17033;
 end   
18'd79804: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=12;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd79805: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=41;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd79806: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=4;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd79807: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=96;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd79808: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=62;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd79809: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd79810: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=51;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd79811: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd79812: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd79813: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16436;
 end   
18'd79814: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16436;
 end   
18'd79815: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16436;
 end   
18'd79816: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16436;
 end   
18'd79817: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16436;
 end   
18'd79818: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16436;
 end   
18'd79942: begin  
rid<=1;
end
18'd79943: begin  
end
18'd79944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd79945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd79946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd79947: begin  
rid<=0;
end
18'd80001: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=45;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3989;
 end   
18'd80002: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=28;
   mapp<=38;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5402;
 end   
18'd80003: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=94;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=7118;
 end   
18'd80004: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=26;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=4684;
 end   
18'd80005: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=78;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd80006: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd80007: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd80142: begin  
rid<=1;
end
18'd80143: begin  
end
18'd80144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd80145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd80146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd80147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd80148: begin  
rid<=0;
end
18'd80201: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=99;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7793;
 end   
18'd80202: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=27;
   mapp<=49;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8856;
 end   
18'd80203: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=92;
   mapp<=57;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9063;
 end   
18'd80204: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=53;
   mapp<=12;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=8197;
 end   
18'd80205: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=95;
   mapp<=1;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=7056;
 end   
18'd80206: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=42;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=7303;
 end   
18'd80207: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=67;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd80208: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=49;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd80209: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=76;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd80210: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=55;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd80211: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd80212: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd80213: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7793;
 end   
18'd80214: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7793;
 end   
18'd80215: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7793;
 end   
18'd80342: begin  
rid<=1;
end
18'd80343: begin  
end
18'd80344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd80345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd80346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd80347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd80348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd80349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd80350: begin  
rid<=0;
end
18'd80401: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=47;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1236;
 end   
18'd80402: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=73;
   mapp<=15;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1204;
 end   
18'd80403: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=65;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=950;
 end   
18'd80404: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=49;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=732;
 end   
18'd80405: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=37;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=1186;
 end   
18'd80406: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=69;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=722;
 end   
18'd80407: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=31;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd80408: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd80409: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd80542: begin  
rid<=1;
end
18'd80543: begin  
end
18'd80544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd80545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd80546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd80547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd80548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd80549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd80550: begin  
rid<=0;
end
18'd80601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=29;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=25639;
 end   
18'd80602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=31;
   mapp<=52;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=25677;
 end   
18'd80603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=78;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd80604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=59;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd80605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=52;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd80606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=89;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd80607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd80608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd80609: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd80610: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd80611: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd80612: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd80613: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25639;
 end   
18'd80742: begin  
rid<=1;
end
18'd80743: begin  
end
18'd80744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd80745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd80746: begin  
rid<=0;
end
18'd80801: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=71;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7858;
 end   
18'd80802: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=47;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6996;
 end   
18'd80803: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=3;
   mapp<=8;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=2630;
 end   
18'd80804: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=11;
   mapp<=56;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=6496;
 end   
18'd80805: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=74;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=5740;
 end   
18'd80806: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=19;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=7164;
 end   
18'd80807: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=7;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=6518;
 end   
18'd80808: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=5;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd80809: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=99;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd80810: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd80811: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd80812: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd80813: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7858;
 end   
18'd80814: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7858;
 end   
18'd80942: begin  
rid<=1;
end
18'd80943: begin  
end
18'd80944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd80945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd80946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd80947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd80948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd80949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd80950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd80951: begin  
rid<=0;
end
18'd81001: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=99;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12514;
 end   
18'd81002: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=54;
   mapp<=92;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=18727;
 end   
18'd81003: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=67;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd81004: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=12;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd81005: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=14;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd81006: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=29;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd81007: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd81008: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd81009: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd81010: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd81011: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd81012: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd81013: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12514;
 end   
18'd81142: begin  
rid<=1;
end
18'd81143: begin  
end
18'd81144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd81145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd81146: begin  
rid<=0;
end
18'd81201: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=74;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=30473;
 end   
18'd81202: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=36;
   mapp<=12;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=24922;
 end   
18'd81203: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=12;
   mapp<=31;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=15240;
 end   
18'd81204: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=87;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd81205: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=57;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd81206: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=3;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd81207: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=91;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd81208: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=82;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd81209: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=29;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd81210: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=27;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd81211: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd81212: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd81213: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=30473;
 end   
18'd81214: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=30473;
 end   
18'd81215: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=30473;
 end   
18'd81216: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=30473;
 end   
18'd81217: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=30473;
 end   
18'd81218: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=30473;
 end   
18'd81342: begin  
rid<=1;
end
18'd81343: begin  
end
18'd81344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd81345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd81346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd81347: begin  
rid<=0;
end
18'd81401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=76;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=26690;
 end   
18'd81402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=24;
   mapp<=46;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=21220;
 end   
18'd81403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=81;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd81404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=95;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd81405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=23;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd81406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=32;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd81407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=43;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd81408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd81409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd81410: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd81411: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd81412: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd81413: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26690;
 end   
18'd81414: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26690;
 end   
18'd81415: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26690;
 end   
18'd81542: begin  
rid<=1;
end
18'd81543: begin  
end
18'd81544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd81545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd81546: begin  
rid<=0;
end
18'd81601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=50;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8613;
 end   
18'd81602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=32;
   mapp<=89;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10099;
 end   
18'd81603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=45;
   mapp<=37;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6613;
 end   
18'd81604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=99;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=9655;
 end   
18'd81605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=35;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=6748;
 end   
18'd81606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=79;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=8068;
 end   
18'd81607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=54;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=8879;
 end   
18'd81608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd81609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd81610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd81611: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd81612: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd81742: begin  
rid<=1;
end
18'd81743: begin  
end
18'd81744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd81745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd81746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd81747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd81748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd81749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd81750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd81751: begin  
rid<=0;
end
18'd81801: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=77;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4299;
 end   
18'd81802: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=5;
   mapp<=90;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2165;
 end   
18'd81803: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=19;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd81804: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=50;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd81805: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd81806: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd81807: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd81942: begin  
rid<=1;
end
18'd81943: begin  
end
18'd81944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd81945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd81946: begin  
rid<=0;
end
18'd82001: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=84;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15194;
 end   
18'd82002: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=51;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11099;
 end   
18'd82003: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=84;
   mapp<=85;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12245;
 end   
18'd82004: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=37;
   mapp<=74;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=15423;
 end   
18'd82005: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=15;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=18783;
 end   
18'd82006: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=89;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=18172;
 end   
18'd82007: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=81;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=15589;
 end   
18'd82008: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=74;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=13364;
 end   
18'd82009: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=59;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd82010: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=50;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd82011: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=46;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd82012: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd82013: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15194;
 end   
18'd82014: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15194;
 end   
18'd82015: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15194;
 end   
18'd82142: begin  
rid<=1;
end
18'd82143: begin  
end
18'd82144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd82145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd82146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd82147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd82148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd82149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd82150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd82151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd82152: begin  
rid<=0;
end
18'd82201: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=21;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=693;
 end   
18'd82202: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=61;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2023;
 end   
18'd82203: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=18;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=614;
 end   
18'd82204: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=46;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=1548;
 end   
18'd82205: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd82342: begin  
rid<=1;
end
18'd82343: begin  
end
18'd82344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd82345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd82346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd82347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd82348: begin  
rid<=0;
end
18'd82401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=60;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3660;
 end   
18'd82402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=46;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=2770;
 end   
18'd82403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=58;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=3500;
 end   
18'd82404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=94;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=5670;
 end   
18'd82405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=71;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=4300;
 end   
18'd82406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=45;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=2750;
 end   
18'd82407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=2;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=180;
 end   
18'd82408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=46;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=2830;
 end   
18'd82409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=20;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=1280;
 end   
18'd82410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=54;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[9]<=3330;
 end   
18'd82411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=53;
   pp<=100;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[10]<=3280;
 end   
18'd82412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd82542: begin  
rid<=1;
end
18'd82543: begin  
end
18'd82544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd82545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd82546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd82547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd82548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd82549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd82550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd82551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd82552: begin  
check<=expctdoutput[8]-outcheck;
end
18'd82553: begin  
check<=expctdoutput[9]-outcheck;
end
18'd82554: begin  
check<=expctdoutput[10]-outcheck;
end
18'd82555: begin  
rid<=0;
end
18'd82601: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=16;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=560;
 end   
18'd82602: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=13;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=465;
 end   
18'd82603: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=35;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1245;
 end   
18'd82604: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=92;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=3250;
 end   
18'd82605: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=18;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=670;
 end   
18'd82606: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=65;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=2325;
 end   
18'd82607: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=70;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=2510;
 end   
18'd82608: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=36;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=1330;
 end   
18'd82609: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=25;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=955;
 end   
18'd82610: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=46;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[9]<=1700;
 end   
18'd82611: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd82742: begin  
rid<=1;
end
18'd82743: begin  
end
18'd82744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd82745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd82746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd82747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd82748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd82749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd82750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd82751: begin  
check<=expctdoutput[7]-outcheck;
end
18'd82752: begin  
check<=expctdoutput[8]-outcheck;
end
18'd82753: begin  
check<=expctdoutput[9]-outcheck;
end
18'd82754: begin  
rid<=0;
end
18'd82801: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=15;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1230;
 end   
18'd82802: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=5;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=420;
 end   
18'd82803: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=26;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=2152;
 end   
18'd82804: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=1;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=112;
 end   
18'd82805: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=73;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=6026;
 end   
18'd82806: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=6;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=542;
 end   
18'd82807: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=80;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=6620;
 end   
18'd82808: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=93;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=7696;
 end   
18'd82809: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=90;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=7460;
 end   
18'd82810: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=91;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[9]<=7552;
 end   
18'd82811: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd82942: begin  
rid<=1;
end
18'd82943: begin  
end
18'd82944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd82945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd82946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd82947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd82948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd82949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd82950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd82951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd82952: begin  
check<=expctdoutput[8]-outcheck;
end
18'd82953: begin  
check<=expctdoutput[9]-outcheck;
end
18'd82954: begin  
rid<=0;
end
18'd83001: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=85;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4845;
 end   
18'd83002: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=10;
 end   
18'd83003: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=49;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=4185;
 end   
18'd83004: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=22;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=1900;
 end   
18'd83005: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd83142: begin  
rid<=1;
end
18'd83143: begin  
end
18'd83144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd83145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd83146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd83147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd83148: begin  
rid<=0;
end
18'd83201: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=92;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=22206;
 end   
18'd83202: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=74;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=23572;
 end   
18'd83203: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=43;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd83204: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=19;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd83205: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=81;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd83206: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=70;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd83207: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=91;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd83208: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=45;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd83209: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd83210: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd83211: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd83212: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd83213: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22206;
 end   
18'd83214: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22206;
 end   
18'd83215: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22206;
 end   
18'd83216: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22206;
 end   
18'd83217: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22206;
 end   
18'd83342: begin  
rid<=1;
end
18'd83343: begin  
end
18'd83344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd83345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd83346: begin  
rid<=0;
end
18'd83401: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=16;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=30319;
 end   
18'd83402: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=8;
   mapp<=79;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=32082;
 end   
18'd83403: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=88;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd83404: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=99;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd83405: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=25;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd83406: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=96;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd83407: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=69;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd83408: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=31;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd83409: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=14;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd83410: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=2;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd83411: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd83412: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd83413: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=30319;
 end   
18'd83414: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=30319;
 end   
18'd83415: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=30319;
 end   
18'd83416: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=30319;
 end   
18'd83417: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=30319;
 end   
18'd83418: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=30319;
 end   
18'd83419: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=30319;
 end   
18'd83542: begin  
rid<=1;
end
18'd83543: begin  
end
18'd83544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd83545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd83546: begin  
rid<=0;
end
18'd83601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=67;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11340;
 end   
18'd83602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=62;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11245;
 end   
18'd83603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=98;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=9748;
 end   
18'd83604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=51;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=8903;
 end   
18'd83605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=88;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=9842;
 end   
18'd83606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=63;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=7557;
 end   
18'd83607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=53;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=3921;
 end   
18'd83608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=5;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=2947;
 end   
18'd83609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd83610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd83611: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd83742: begin  
rid<=1;
end
18'd83743: begin  
end
18'd83744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd83745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd83746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd83747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd83748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd83749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd83750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd83751: begin  
check<=expctdoutput[7]-outcheck;
end
18'd83752: begin  
rid<=0;
end
18'd83801: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=18;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2340;
 end   
18'd83802: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=35;
   mapp<=18;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2854;
 end   
18'd83803: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=72;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=4606;
 end   
18'd83804: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=94;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=4172;
 end   
18'd83805: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=70;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=2630;
 end   
18'd83806: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=38;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=1469;
 end   
18'd83807: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=21;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=2013;
 end   
18'd83808: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=45;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=1685;
 end   
18'd83809: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=23;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=1999;
 end   
18'd83810: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=43;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[9]<=3139;
 end   
18'd83811: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd83812: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd83813: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=2340;
 end   
18'd83942: begin  
rid<=1;
end
18'd83943: begin  
end
18'd83944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd83945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd83946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd83947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd83948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd83949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd83950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd83951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd83952: begin  
check<=expctdoutput[8]-outcheck;
end
18'd83953: begin  
check<=expctdoutput[9]-outcheck;
end
18'd83954: begin  
rid<=0;
end
18'd84001: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=18;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8682;
 end   
18'd84002: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=75;
   mapp<=92;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5716;
 end   
18'd84003: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=54;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=2792;
 end   
18'd84004: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=24;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=2787;
 end   
18'd84005: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=31;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=5548;
 end   
18'd84006: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=66;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=3413;
 end   
18'd84007: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=29;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=2232;
 end   
18'd84008: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=22;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=4666;
 end   
18'd84009: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd84010: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd84011: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd84142: begin  
rid<=1;
end
18'd84143: begin  
end
18'd84144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd84145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd84146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd84147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd84148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd84149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd84150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd84151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd84152: begin  
rid<=0;
end
18'd84201: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=38;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11068;
 end   
18'd84202: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=75;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10988;
 end   
18'd84203: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=44;
   mapp<=28;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=11957;
 end   
18'd84204: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=25;
   mapp<=22;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=15169;
 end   
18'd84205: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=39;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd84206: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=21;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd84207: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=40;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd84208: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd84209: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd84210: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd84211: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd84212: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd84213: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11068;
 end   
18'd84214: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11068;
 end   
18'd84215: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11068;
 end   
18'd84216: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11068;
 end   
18'd84217: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11068;
 end   
18'd84342: begin  
rid<=1;
end
18'd84343: begin  
end
18'd84344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd84345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd84346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd84347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd84348: begin  
rid<=0;
end
18'd84401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=76;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9157;
 end   
18'd84402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=40;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6711;
 end   
18'd84403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=23;
   mapp<=47;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5793;
 end   
18'd84404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=51;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=5359;
 end   
18'd84405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=7;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=2842;
 end   
18'd84406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=51;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=5637;
 end   
18'd84407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=10;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=4871;
 end   
18'd84408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=57;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=7689;
 end   
18'd84409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=77;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=6361;
 end   
18'd84410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd84411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd84412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd84413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9157;
 end   
18'd84414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9157;
 end   
18'd84542: begin  
rid<=1;
end
18'd84543: begin  
end
18'd84544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd84545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd84546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd84547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd84548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd84549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd84550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd84551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd84552: begin  
check<=expctdoutput[8]-outcheck;
end
18'd84553: begin  
rid<=0;
end
18'd84601: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=99;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9669;
 end   
18'd84602: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=48;
   mapp<=6;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9707;
 end   
18'd84603: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=30;
   mapp<=85;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=7458;
 end   
18'd84604: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=73;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=6775;
 end   
18'd84605: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=58;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=11278;
 end   
18'd84606: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=16;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=7863;
 end   
18'd84607: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=84;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=8929;
 end   
18'd84608: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=73;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=5633;
 end   
18'd84609: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=31;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=9298;
 end   
18'd84610: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=4;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd84611: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=83;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd84612: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd84613: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9669;
 end   
18'd84614: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9669;
 end   
18'd84742: begin  
rid<=1;
end
18'd84743: begin  
end
18'd84744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd84745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd84746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd84747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd84748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd84749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd84750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd84751: begin  
check<=expctdoutput[7]-outcheck;
end
18'd84752: begin  
check<=expctdoutput[8]-outcheck;
end
18'd84753: begin  
rid<=0;
end
18'd84801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=9;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5049;
 end   
18'd84802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=57;
   mapp<=87;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4441;
 end   
18'd84803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=64;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=4472;
 end   
18'd84804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=68;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=6000;
 end   
18'd84805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=94;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=5389;
 end   
18'd84806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=79;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=2072;
 end   
18'd84807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd84808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd84809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd84942: begin  
rid<=1;
end
18'd84943: begin  
end
18'd84944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd84945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd84946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd84947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd84948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd84949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd84950: begin  
rid<=0;
end
18'd85001: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=17;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6488;
 end   
18'd85002: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=9;
   mapp<=23;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4598;
 end   
18'd85003: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=43;
   mapp<=72;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6284;
 end   
18'd85004: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=67;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd85005: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd85006: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd85007: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd85008: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd85009: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd85010: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd85142: begin  
rid<=1;
end
18'd85143: begin  
end
18'd85144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd85145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd85146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd85147: begin  
rid<=0;
end
18'd85201: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=69;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6279;
 end   
18'd85202: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=38;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3468;
 end   
18'd85203: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=4;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=384;
 end   
18'd85204: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=76;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=6946;
 end   
18'd85205: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=12;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=1132;
 end   
18'd85206: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=91;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=8331;
 end   
18'd85207: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=93;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=8523;
 end   
18'd85208: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=9;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=889;
 end   
18'd85209: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=20;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=1900;
 end   
18'd85210: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd85342: begin  
rid<=1;
end
18'd85343: begin  
end
18'd85344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd85345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd85346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd85347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd85348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd85349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd85350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd85351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd85352: begin  
check<=expctdoutput[8]-outcheck;
end
18'd85353: begin  
rid<=0;
end
18'd85401: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=89;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4970;
 end   
18'd85402: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=94;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7320;
 end   
18'd85403: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=42;
   mapp<=59;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=10899;
 end   
18'd85404: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd85405: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd85406: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd85407: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd85408: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd85542: begin  
rid<=1;
end
18'd85543: begin  
end
18'd85544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd85545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd85546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd85547: begin  
rid<=0;
end
18'd85601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=45;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13833;
 end   
18'd85602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=88;
   mapp<=64;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=15098;
 end   
18'd85603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=49;
   mapp<=86;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=14027;
 end   
18'd85604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=27;
   mapp<=71;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=12241;
 end   
18'd85605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd85606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd85607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd85608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd85609: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd85610: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd85611: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd85742: begin  
rid<=1;
end
18'd85743: begin  
end
18'd85744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd85745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd85746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd85747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd85748: begin  
rid<=0;
end
18'd85801: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=46;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3726;
 end   
18'd85802: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd85942: begin  
rid<=1;
end
18'd85943: begin  
end
18'd85944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd85945: begin  
rid<=0;
end
18'd86001: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=68;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13596;
 end   
18'd86002: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=89;
   mapp<=50;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=16788;
 end   
18'd86003: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=83;
   mapp<=32;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=23039;
 end   
18'd86004: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=9;
   mapp<=73;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=21031;
 end   
18'd86005: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=87;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd86006: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=95;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd86007: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd86008: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd86009: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd86010: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd86011: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd86012: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd86013: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13596;
 end   
18'd86014: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13596;
 end   
18'd86015: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13596;
 end   
18'd86142: begin  
rid<=1;
end
18'd86143: begin  
end
18'd86144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd86145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd86146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd86147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd86148: begin  
rid<=0;
end
18'd86201: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=48;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4637;
 end   
18'd86202: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=79;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3336;
 end   
18'd86203: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=7;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1343;
 end   
18'd86204: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=30;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=3090;
 end   
18'd86205: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=54;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=2181;
 end   
18'd86206: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=1;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=1489;
 end   
18'd86207: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=40;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=3125;
 end   
18'd86208: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=43;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=2377;
 end   
18'd86209: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=18;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=1202;
 end   
18'd86210: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd86211: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd86212: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd86342: begin  
rid<=1;
end
18'd86343: begin  
end
18'd86344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd86345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd86346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd86347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd86348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd86349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd86350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd86351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd86352: begin  
check<=expctdoutput[8]-outcheck;
end
18'd86353: begin  
rid<=0;
end
18'd86401: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=83;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5976;
 end   
18'd86402: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=85;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6130;
 end   
18'd86403: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=86;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6212;
 end   
18'd86404: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=20;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=1470;
 end   
18'd86405: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd86542: begin  
rid<=1;
end
18'd86543: begin  
end
18'd86544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd86545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd86546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd86547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd86548: begin  
rid<=0;
end
18'd86601: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=6;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15374;
 end   
18'd86602: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=21;
   mapp<=6;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=14814;
 end   
18'd86603: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=75;
   mapp<=76;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=16027;
 end   
18'd86604: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=20;
   mapp<=24;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=19119;
 end   
18'd86605: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=92;
   mapp<=52;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=16205;
 end   
18'd86606: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=65;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd86607: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=47;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd86608: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd86609: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd86610: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd86611: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd86612: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd86613: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15374;
 end   
18'd86614: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15374;
 end   
18'd86615: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15374;
 end   
18'd86616: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15374;
 end   
18'd86617: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15374;
 end   
18'd86618: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15374;
 end   
18'd86742: begin  
rid<=1;
end
18'd86743: begin  
end
18'd86744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd86745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd86746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd86747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd86748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd86749: begin  
rid<=0;
end
18'd86801: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=62;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6739;
 end   
18'd86802: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=89;
   mapp<=29;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9386;
 end   
18'd86803: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=23;
   mapp<=82;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6617;
 end   
18'd86804: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=70;
   mapp<=5;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=10622;
 end   
18'd86805: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=42;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=11992;
 end   
18'd86806: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=82;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=12281;
 end   
18'd86807: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=96;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd86808: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=80;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd86809: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=69;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd86810: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd86811: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd86812: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd86813: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6739;
 end   
18'd86942: begin  
rid<=1;
end
18'd86943: begin  
end
18'd86944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd86945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd86946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd86947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd86948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd86949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd86950: begin  
rid<=0;
end
18'd87001: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=37;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12020;
 end   
18'd87002: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=1;
   mapp<=36;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11271;
 end   
18'd87003: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=76;
   mapp<=55;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=10314;
 end   
18'd87004: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=4;
   mapp<=74;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=13051;
 end   
18'd87005: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=73;
   mapp<=77;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=9198;
 end   
18'd87006: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=54;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=13550;
 end   
18'd87007: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd87008: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd87009: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd87010: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd87011: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd87012: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd87013: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12020;
 end   
18'd87014: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12020;
 end   
18'd87015: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12020;
 end   
18'd87142: begin  
rid<=1;
end
18'd87143: begin  
end
18'd87144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd87145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd87146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd87147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd87148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd87149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd87150: begin  
rid<=0;
end
18'd87201: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=18;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1710;
 end   
18'd87202: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=25;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=460;
 end   
18'd87203: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=85;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=1550;
 end   
18'd87204: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=62;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=1146;
 end   
18'd87205: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=29;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=562;
 end   
18'd87206: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=60;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=1130;
 end   
18'd87207: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd87342: begin  
rid<=1;
end
18'd87343: begin  
end
18'd87344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd87345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd87346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd87347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd87348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd87349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd87350: begin  
rid<=0;
end
18'd87401: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=62;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=558;
 end   
18'd87402: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=24;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=226;
 end   
18'd87403: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=74;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=686;
 end   
18'd87404: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=82;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=768;
 end   
18'd87405: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=75;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=715;
 end   
18'd87406: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=15;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=185;
 end   
18'd87407: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd87542: begin  
rid<=1;
end
18'd87543: begin  
end
18'd87544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd87545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd87546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd87547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd87548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd87549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd87550: begin  
rid<=0;
end
18'd87601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=89;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6316;
 end   
18'd87602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=51;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10346;
 end   
18'd87603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=84;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=10607;
 end   
18'd87604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=61;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=9131;
 end   
18'd87605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=72;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=10834;
 end   
18'd87606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=86;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=11070;
 end   
18'd87607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd87608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd87609: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd87742: begin  
rid<=1;
end
18'd87743: begin  
end
18'd87744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd87745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd87746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd87747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd87748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd87749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd87750: begin  
rid<=0;
end
18'd87801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=17;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=22924;
 end   
18'd87802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=64;
   mapp<=76;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=21042;
 end   
18'd87803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=16;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd87804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=14;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd87805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=66;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd87806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=96;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd87807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=73;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd87808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=48;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd87809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd87810: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd87811: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd87812: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd87813: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22924;
 end   
18'd87814: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22924;
 end   
18'd87815: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22924;
 end   
18'd87942: begin  
rid<=1;
end
18'd87943: begin  
end
18'd87944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd87945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd87946: begin  
rid<=0;
end
18'd88001: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=89;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5469;
 end   
18'd88002: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=20;
   mapp<=91;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9429;
 end   
18'd88003: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd88004: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd88005: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd88142: begin  
rid<=1;
end
18'd88143: begin  
end
18'd88144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd88145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd88146: begin  
rid<=0;
end
18'd88201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=25;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8726;
 end   
18'd88202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=28;
   mapp<=81;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11185;
 end   
18'd88203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=73;
   mapp<=71;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8756;
 end   
18'd88204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=54;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=5643;
 end   
18'd88205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=9;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=5627;
 end   
18'd88206: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=30;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=11119;
 end   
18'd88207: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=38;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=12138;
 end   
18'd88208: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=91;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=11633;
 end   
18'd88209: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=39;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd88210: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=53;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd88211: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd88212: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd88213: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8726;
 end   
18'd88342: begin  
rid<=1;
end
18'd88343: begin  
end
18'd88344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd88345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd88346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd88347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd88348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd88349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd88350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd88351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd88352: begin  
rid<=0;
end
18'd88401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=39;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=24340;
 end   
18'd88402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=85;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=25192;
 end   
18'd88403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=41;
   mapp<=90;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=24462;
 end   
18'd88404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=67;
   mapp<=97;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=20929;
 end   
18'd88405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=20;
   mapp<=56;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=18692;
 end   
18'd88406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=60;
   mapp<=73;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=21276;
 end   
18'd88407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd88408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd88409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd88410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd88411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd88412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd88413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24340;
 end   
18'd88414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24340;
 end   
18'd88415: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24340;
 end   
18'd88416: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24340;
 end   
18'd88417: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24340;
 end   
18'd88542: begin  
rid<=1;
end
18'd88543: begin  
end
18'd88544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd88545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd88546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd88547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd88548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd88549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd88550: begin  
rid<=0;
end
18'd88601: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=60;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15997;
 end   
18'd88602: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=62;
   mapp<=6;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=17275;
 end   
18'd88603: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=32;
   mapp<=89;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12384;
 end   
18'd88604: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=92;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd88605: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=43;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd88606: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=63;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd88607: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd88608: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd88609: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd88610: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd88611: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd88612: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd88742: begin  
rid<=1;
end
18'd88743: begin  
end
18'd88744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd88745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd88746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd88747: begin  
rid<=0;
end
18'd88801: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=49;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5024;
 end   
18'd88802: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=12;
   mapp<=43;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2957;
 end   
18'd88803: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=3678;
 end   
18'd88804: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd88805: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd88806: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd88942: begin  
rid<=1;
end
18'd88943: begin  
end
18'd88944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd88945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd88946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd88947: begin  
rid<=0;
end
18'd89001: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=38;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=17879;
 end   
18'd89002: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=23;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=12369;
 end   
18'd89003: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=5;
   mapp<=3;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=7955;
 end   
18'd89004: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=11;
   mapp<=64;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=18765;
 end   
18'd89005: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=93;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd89006: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=17;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd89007: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=43;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd89008: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=27;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd89009: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=14;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd89010: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=90;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd89011: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd89012: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd89013: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17879;
 end   
18'd89014: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17879;
 end   
18'd89015: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17879;
 end   
18'd89016: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17879;
 end   
18'd89017: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17879;
 end   
18'd89142: begin  
rid<=1;
end
18'd89143: begin  
end
18'd89144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd89145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd89146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd89147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd89148: begin  
rid<=0;
end
18'd89201: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=44;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1716;
 end   
18'd89202: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd89342: begin  
rid<=1;
end
18'd89343: begin  
end
18'd89344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd89345: begin  
rid<=0;
end
18'd89401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=37;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7011;
 end   
18'd89402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=34;
   mapp<=33;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8561;
 end   
18'd89403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=77;
   mapp<=40;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=10410;
 end   
18'd89404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=71;
   mapp<=1;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=7572;
 end   
18'd89405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=83;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=8800;
 end   
18'd89406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd89407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd89408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd89409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd89410: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd89411: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd89412: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd89542: begin  
rid<=1;
end
18'd89543: begin  
end
18'd89544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd89545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd89546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd89547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd89548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd89549: begin  
rid<=0;
end
18'd89601: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=5;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11489;
 end   
18'd89602: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=1;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10686;
 end   
18'd89603: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=34;
   mapp<=68;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=11833;
 end   
18'd89604: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=70;
   mapp<=82;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=10923;
 end   
18'd89605: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=55;
   mapp<=48;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=8983;
 end   
18'd89606: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=7;
   mapp<=66;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=9395;
 end   
18'd89607: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd89608: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd89609: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd89610: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd89611: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd89612: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd89613: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11489;
 end   
18'd89614: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11489;
 end   
18'd89615: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11489;
 end   
18'd89616: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11489;
 end   
18'd89617: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11489;
 end   
18'd89742: begin  
rid<=1;
end
18'd89743: begin  
end
18'd89744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd89745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd89746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd89747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd89748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd89749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd89750: begin  
rid<=0;
end
18'd89801: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=87;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=26596;
 end   
18'd89802: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=64;
   mapp<=3;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=21463;
 end   
18'd89803: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=13;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd89804: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=13;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd89805: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=52;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd89806: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=70;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd89807: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=78;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd89808: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=66;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd89809: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=4;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd89810: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd89811: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd89812: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd89813: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26596;
 end   
18'd89814: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26596;
 end   
18'd89815: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26596;
 end   
18'd89816: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26596;
 end   
18'd89817: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26596;
 end   
18'd89818: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26596;
 end   
18'd89819: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26596;
 end   
18'd89942: begin  
rid<=1;
end
18'd89943: begin  
end
18'd89944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd89945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd89946: begin  
rid<=0;
end
18'd90001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=55;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=20340;
 end   
18'd90002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=90;
   mapp<=37;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13103;
 end   
18'd90003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=46;
   mapp<=37;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=15940;
 end   
18'd90004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=82;
   mapp<=59;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=13446;
 end   
18'd90005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=35;
   mapp<=32;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=16545;
 end   
18'd90006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=93;
   mapp<=55;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=11367;
 end   
18'd90007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd90008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd90009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd90010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd90011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd90012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd90013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20340;
 end   
18'd90014: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20340;
 end   
18'd90015: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20340;
 end   
18'd90016: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20340;
 end   
18'd90017: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20340;
 end   
18'd90142: begin  
rid<=1;
end
18'd90143: begin  
end
18'd90144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd90145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd90146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd90147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd90148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd90149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd90150: begin  
rid<=0;
end
18'd90201: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=63;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12667;
 end   
18'd90202: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=49;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=18845;
 end   
18'd90203: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=76;
   mapp<=3;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=17348;
 end   
18'd90204: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=97;
   mapp<=14;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=16092;
 end   
18'd90205: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=34;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd90206: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=47;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd90207: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=26;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd90208: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd90209: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd90210: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd90211: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd90212: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd90213: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12667;
 end   
18'd90214: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12667;
 end   
18'd90215: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12667;
 end   
18'd90216: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12667;
 end   
18'd90217: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12667;
 end   
18'd90342: begin  
rid<=1;
end
18'd90343: begin  
end
18'd90344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd90345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd90346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd90347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd90348: begin  
rid<=0;
end
18'd90401: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=69;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10923;
 end   
18'd90402: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=75;
   mapp<=61;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9289;
 end   
18'd90403: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=39;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9464;
 end   
18'd90404: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=96;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=13803;
 end   
18'd90405: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=81;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=11823;
 end   
18'd90406: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=71;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=10730;
 end   
18'd90407: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=68;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=7109;
 end   
18'd90408: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=13;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=5292;
 end   
18'd90409: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=66;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=7982;
 end   
18'd90410: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=30;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[9]<=3216;
 end   
18'd90411: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=6;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd90412: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd90413: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10923;
 end   
18'd90542: begin  
rid<=1;
end
18'd90543: begin  
end
18'd90544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd90545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd90546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd90547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd90548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd90549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd90550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd90551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd90552: begin  
check<=expctdoutput[8]-outcheck;
end
18'd90553: begin  
check<=expctdoutput[9]-outcheck;
end
18'd90554: begin  
rid<=0;
end
18'd90601: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=91;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=17597;
 end   
18'd90602: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=93;
   mapp<=84;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=17596;
 end   
18'd90603: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=96;
   mapp<=46;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9981;
 end   
18'd90604: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=59;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=6254;
 end   
18'd90605: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd90606: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd90607: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd90608: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd90609: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd90742: begin  
rid<=1;
end
18'd90743: begin  
end
18'd90744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd90745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd90746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd90747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd90748: begin  
rid<=0;
end
18'd90801: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=67;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7014;
 end   
18'd90802: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=69;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6254;
 end   
18'd90803: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=65;
   mapp<=12;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=4706;
 end   
18'd90804: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=3;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=3848;
 end   
18'd90805: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=73;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=7578;
 end   
18'd90806: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=91;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=6385;
 end   
18'd90807: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=16;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=2867;
 end   
18'd90808: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=49;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=3604;
 end   
18'd90809: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=15;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd90810: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=18;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd90811: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd90812: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd90813: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7014;
 end   
18'd90942: begin  
rid<=1;
end
18'd90943: begin  
end
18'd90944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd90945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd90946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd90947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd90948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd90949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd90950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd90951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd90952: begin  
rid<=0;
end
18'd91001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=36;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3492;
 end   
18'd91002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=11;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=406;
 end   
18'd91003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=91;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=3296;
 end   
18'd91004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=74;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=2694;
 end   
18'd91005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=63;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=2308;
 end   
18'd91006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=25;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=950;
 end   
18'd91007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=7;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=312;
 end   
18'd91008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=70;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=2590;
 end   
18'd91009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=21;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=836;
 end   
18'd91010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=27;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[9]<=1062;
 end   
18'd91011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=58;
   pp<=100;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[10]<=2188;
 end   
18'd91012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd91142: begin  
rid<=1;
end
18'd91143: begin  
end
18'd91144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd91145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd91146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd91147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd91148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd91149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd91150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd91151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd91152: begin  
check<=expctdoutput[8]-outcheck;
end
18'd91153: begin  
check<=expctdoutput[9]-outcheck;
end
18'd91154: begin  
check<=expctdoutput[10]-outcheck;
end
18'd91155: begin  
rid<=0;
end
18'd91201: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=12;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=912;
 end   
18'd91202: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=99;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=1198;
 end   
18'd91203: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=19;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=248;
 end   
18'd91204: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=41;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=522;
 end   
18'd91205: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=11;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=172;
 end   
18'd91206: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd91342: begin  
rid<=1;
end
18'd91343: begin  
end
18'd91344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd91345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd91346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd91347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd91348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd91349: begin  
rid<=0;
end
18'd91401: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=83;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8825;
 end   
18'd91402: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=32;
   mapp<=30;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5392;
 end   
18'd91403: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=88;
   mapp<=14;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9324;
 end   
18'd91404: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=39;
   mapp<=36;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=5057;
 end   
18'd91405: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=5;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=5463;
 end   
18'd91406: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd91407: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=40;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd91408: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=68;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd91409: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd91410: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd91411: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd91412: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd91542: begin  
rid<=1;
end
18'd91543: begin  
end
18'd91544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd91545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd91546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd91547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd91548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd91549: begin  
rid<=0;
end
18'd91601: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=37;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3145;
 end   
18'd91602: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=20;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1710;
 end   
18'd91603: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=24;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=2060;
 end   
18'd91604: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=97;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=8275;
 end   
18'd91605: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=54;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=4630;
 end   
18'd91606: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=3;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=305;
 end   
18'd91607: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=94;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=8050;
 end   
18'd91608: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd91742: begin  
rid<=1;
end
18'd91743: begin  
end
18'd91744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd91745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd91746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd91747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd91748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd91749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd91750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd91751: begin  
rid<=0;
end
18'd91801: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=94;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6986;
 end   
18'd91802: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=26;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4433;
 end   
18'd91803: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=63;
   mapp<=2;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6103;
 end   
18'd91804: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=28;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd91805: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=48;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd91806: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=79;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd91807: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=51;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd91808: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd91809: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd91810: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd91811: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd91812: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd91942: begin  
rid<=1;
end
18'd91943: begin  
end
18'd91944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd91945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd91946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd91947: begin  
rid<=0;
end
18'd92001: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=98;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14006;
 end   
18'd92002: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=58;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd92003: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=30;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd92004: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=53;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd92005: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd92006: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd92007: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd92008: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd92142: begin  
rid<=1;
end
18'd92143: begin  
end
18'd92144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd92145: begin  
rid<=0;
end
18'd92201: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=58;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=18179;
 end   
18'd92202: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=52;
   mapp<=49;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=16134;
 end   
18'd92203: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=29;
   mapp<=85;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=16746;
 end   
18'd92204: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=40;
   mapp<=55;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=15251;
 end   
18'd92205: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=60;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd92206: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=46;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd92207: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=27;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd92208: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=44;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd92209: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=22;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd92210: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd92211: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd92212: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd92213: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18179;
 end   
18'd92214: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18179;
 end   
18'd92215: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18179;
 end   
18'd92342: begin  
rid<=1;
end
18'd92343: begin  
end
18'd92344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd92345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd92346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd92347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd92348: begin  
rid<=0;
end
18'd92401: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=76;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=17735;
 end   
18'd92402: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=80;
   mapp<=33;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=19511;
 end   
18'd92403: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=69;
   mapp<=56;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=18526;
 end   
18'd92404: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=88;
   mapp<=51;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=16898;
 end   
18'd92405: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=29;
   mapp<=91;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=16042;
 end   
18'd92406: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=34;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=13642;
 end   
18'd92407: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd92408: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd92409: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd92410: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd92411: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd92412: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd92413: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17735;
 end   
18'd92414: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17735;
 end   
18'd92415: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17735;
 end   
18'd92542: begin  
rid<=1;
end
18'd92543: begin  
end
18'd92544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd92545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd92546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd92547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd92548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd92549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd92550: begin  
rid<=0;
end
18'd92601: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=74;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2360;
 end   
18'd92602: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=60;
   mapp<=27;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3283;
 end   
18'd92603: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=99;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd92604: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd92605: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd92742: begin  
rid<=1;
end
18'd92743: begin  
end
18'd92744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd92745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd92746: begin  
rid<=0;
end
18'd92801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=23;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=27826;
 end   
18'd92802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=1;
   mapp<=65;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=26424;
 end   
18'd92803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=87;
   mapp<=28;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=35535;
 end   
18'd92804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=88;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd92805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=97;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd92806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=52;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd92807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=75;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd92808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=50;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd92809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=78;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd92810: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd92811: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd92812: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd92813: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=27826;
 end   
18'd92814: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=27826;
 end   
18'd92815: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=27826;
 end   
18'd92816: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=27826;
 end   
18'd92942: begin  
rid<=1;
end
18'd92943: begin  
end
18'd92944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd92945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd92946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd92947: begin  
rid<=0;
end
18'd93001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=21;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7181;
 end   
18'd93002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=27;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd93003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=64;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd93004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=40;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd93005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=13;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd93006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd93007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd93008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd93009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd93010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd93142: begin  
rid<=1;
end
18'd93143: begin  
end
18'd93144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd93145: begin  
rid<=0;
end
18'd93201: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=22;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13707;
 end   
18'd93202: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=16;
   mapp<=63;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10918;
 end   
18'd93203: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=54;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd93204: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=86;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd93205: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=25;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd93206: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=24;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd93207: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=18;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd93208: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd93209: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd93210: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd93211: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd93212: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd93213: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13707;
 end   
18'd93214: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13707;
 end   
18'd93215: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13707;
 end   
18'd93342: begin  
rid<=1;
end
18'd93343: begin  
end
18'd93344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd93345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd93346: begin  
rid<=0;
end
18'd93401: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=88;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5192;
 end   
18'd93402: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=82;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4848;
 end   
18'd93403: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=41;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=2439;
 end   
18'd93404: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd93542: begin  
rid<=1;
end
18'd93543: begin  
end
18'd93544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd93545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd93546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd93547: begin  
rid<=0;
end
18'd93601: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=22;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1452;
 end   
18'd93602: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=54;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3574;
 end   
18'd93603: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=52;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=3452;
 end   
18'd93604: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=50;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=3330;
 end   
18'd93605: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=16;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=1096;
 end   
18'd93606: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=26;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=1766;
 end   
18'd93607: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=86;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=5736;
 end   
18'd93608: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=2;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=202;
 end   
18'd93609: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=37;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=2522;
 end   
18'd93610: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=1;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[9]<=156;
 end   
18'd93611: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=1;
   mapp<=0;
   pp<=100;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[10]<=166;
 end   
18'd93612: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd93742: begin  
rid<=1;
end
18'd93743: begin  
end
18'd93744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd93745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd93746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd93747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd93748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd93749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd93750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd93751: begin  
check<=expctdoutput[7]-outcheck;
end
18'd93752: begin  
check<=expctdoutput[8]-outcheck;
end
18'd93753: begin  
check<=expctdoutput[9]-outcheck;
end
18'd93754: begin  
check<=expctdoutput[10]-outcheck;
end
18'd93755: begin  
rid<=0;
end
18'd93801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=81;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2957;
 end   
18'd93802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=43;
   mapp<=65;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=746;
 end   
18'd93803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=10;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=560;
 end   
18'd93804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=8;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=5831;
 end   
18'd93805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=89;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=3988;
 end   
18'd93806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=58;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=5626;
 end   
18'd93807: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=84;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd93808: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd93809: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd93942: begin  
rid<=1;
end
18'd93943: begin  
end
18'd93944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd93945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd93946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd93947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd93948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd93949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd93950: begin  
rid<=0;
end
18'd94001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=18;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=23416;
 end   
18'd94002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=73;
   mapp<=87;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=29142;
 end   
18'd94003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=53;
   mapp<=71;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=25603;
 end   
18'd94004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=81;
   mapp<=90;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=24048;
 end   
18'd94005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=62;
   mapp<=72;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=20317;
 end   
18'd94006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=96;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd94007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=13;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd94008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=51;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd94009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=15;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd94010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd94011: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd94012: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd94013: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23416;
 end   
18'd94014: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23416;
 end   
18'd94142: begin  
rid<=1;
end
18'd94143: begin  
end
18'd94144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd94145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd94146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd94147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd94148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd94149: begin  
rid<=0;
end
18'd94201: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=84;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8281;
 end   
18'd94202: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=33;
   mapp<=64;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11129;
 end   
18'd94203: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=72;
   mapp<=4;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9527;
 end   
18'd94204: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=21;
   mapp<=37;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=10592;
 end   
18'd94205: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=44;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd94206: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd94207: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=57;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd94208: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd94209: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd94210: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd94211: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd94212: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd94213: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8281;
 end   
18'd94342: begin  
rid<=1;
end
18'd94343: begin  
end
18'd94344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd94345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd94346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd94347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd94348: begin  
rid<=0;
end
18'd94401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=43;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3499;
 end   
18'd94402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=76;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd94403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=31;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd94404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd94405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd94406: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd94542: begin  
rid<=1;
end
18'd94543: begin  
end
18'd94544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd94545: begin  
rid<=0;
end
18'd94601: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=53;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=689;
 end   
18'd94602: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=11;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=153;
 end   
18'd94603: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=93;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1229;
 end   
18'd94604: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=32;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=446;
 end   
18'd94605: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=51;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=703;
 end   
18'd94606: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=14;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=232;
 end   
18'd94607: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=99;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=1347;
 end   
18'd94608: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd94742: begin  
rid<=1;
end
18'd94743: begin  
end
18'd94744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd94745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd94746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd94747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd94748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd94749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd94750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd94751: begin  
rid<=0;
end
18'd94801: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=69;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7285;
 end   
18'd94802: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=35;
   mapp<=49;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5955;
 end   
18'd94803: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=62;
   mapp<=52;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6570;
 end   
18'd94804: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=12;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=2851;
 end   
18'd94805: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=41;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=6284;
 end   
18'd94806: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=9;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=7381;
 end   
18'd94807: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd94808: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd94809: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd94810: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd94811: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd94942: begin  
rid<=1;
end
18'd94943: begin  
end
18'd94944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd94945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd94946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd94947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd94948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd94949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd94950: begin  
rid<=0;
end
18'd95001: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=63;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1302;
 end   
18'd95002: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=21;
   mapp<=11;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=433;
 end   
18'd95003: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=6;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=617;
 end   
18'd95004: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=45;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=1268;
 end   
18'd95005: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=43;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=1321;
 end   
18'd95006: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=50;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=1923;
 end   
18'd95007: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=93;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=2345;
 end   
18'd95008: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=64;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=1620;
 end   
18'd95009: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=42;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=1278;
 end   
18'd95010: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=44;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd95011: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd95012: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd95142: begin  
rid<=1;
end
18'd95143: begin  
end
18'd95144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd95145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd95146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd95147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd95148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd95149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd95150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd95151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd95152: begin  
check<=expctdoutput[8]-outcheck;
end
18'd95153: begin  
rid<=0;
end
18'd95201: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=6;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2798;
 end   
18'd95202: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=43;
   mapp<=25;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4234;
 end   
18'd95203: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=29;
   mapp<=59;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=2856;
 end   
18'd95204: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd95205: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd95206: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd95207: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd95208: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd95342: begin  
rid<=1;
end
18'd95343: begin  
end
18'd95344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd95345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd95346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd95347: begin  
rid<=0;
end
18'd95401: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=41;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5547;
 end   
18'd95402: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=59;
   mapp<=28;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6175;
 end   
18'd95403: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=20;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=2340;
 end   
18'd95404: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=15;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=2687;
 end   
18'd95405: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=44;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=6404;
 end   
18'd95406: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=78;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd95407: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd95408: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd95542: begin  
rid<=1;
end
18'd95543: begin  
end
18'd95544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd95545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd95546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd95547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd95548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd95549: begin  
rid<=0;
end
18'd95601: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=37;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5451;
 end   
18'd95602: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=35;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6946;
 end   
18'd95603: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=30;
   mapp<=38;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8536;
 end   
18'd95604: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=82;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=7431;
 end   
18'd95605: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=15;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd95606: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=80;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd95607: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd95608: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd95609: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd95742: begin  
rid<=1;
end
18'd95743: begin  
end
18'd95744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd95745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd95746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd95747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd95748: begin  
rid<=0;
end
18'd95801: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=94;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10930;
 end   
18'd95802: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=29;
   mapp<=4;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7886;
 end   
18'd95803: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=32;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd95804: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=9;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd95805: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=16;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd95806: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=29;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd95807: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=61;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd95808: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=33;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd95809: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd95810: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd95811: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd95812: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd95813: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10930;
 end   
18'd95814: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10930;
 end   
18'd95815: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10930;
 end   
18'd95816: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10930;
 end   
18'd95817: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10930;
 end   
18'd95942: begin  
rid<=1;
end
18'd95943: begin  
end
18'd95944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd95945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd95946: begin  
rid<=0;
end
18'd96001: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=87;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=21757;
 end   
18'd96002: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=70;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=19169;
 end   
18'd96003: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=89;
   mapp<=73;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=21349;
 end   
18'd96004: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=29;
   mapp<=39;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=20579;
 end   
18'd96005: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=60;
   mapp<=80;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=20835;
 end   
18'd96006: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=21;
   mapp<=35;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=21982;
 end   
18'd96007: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=97;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd96008: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd96009: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=63;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd96010: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=44;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd96011: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=21;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd96012: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd96013: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21757;
 end   
18'd96014: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21757;
 end   
18'd96015: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21757;
 end   
18'd96016: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21757;
 end   
18'd96017: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21757;
 end   
18'd96142: begin  
rid<=1;
end
18'd96143: begin  
end
18'd96144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd96145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd96146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd96147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd96148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd96149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd96150: begin  
rid<=0;
end
18'd96201: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=37;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=26499;
 end   
18'd96202: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=31;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd96203: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=55;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd96204: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=51;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd96205: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=51;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd96206: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=90;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd96207: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=52;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd96208: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=95;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd96209: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=20;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd96210: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=61;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd96211: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=60;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd96212: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd96213: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26499;
 end   
18'd96214: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26499;
 end   
18'd96215: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26499;
 end   
18'd96216: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26499;
 end   
18'd96217: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26499;
 end   
18'd96218: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26499;
 end   
18'd96219: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26499;
 end   
18'd96220: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26499;
 end   
18'd96221: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26499;
 end   
18'd96222: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26499;
 end   
18'd96342: begin  
rid<=1;
end
18'd96343: begin  
end
18'd96344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd96345: begin  
rid<=0;
end
18'd96401: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=91;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3127;
 end   
18'd96402: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=1;
   mapp<=33;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2618;
 end   
18'd96403: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=78;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5543;
 end   
18'd96404: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=87;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=5595;
 end   
18'd96405: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=79;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=2726;
 end   
18'd96406: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd96407: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd96408: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd96542: begin  
rid<=1;
end
18'd96543: begin  
end
18'd96544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd96545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd96546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd96547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd96548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd96549: begin  
rid<=0;
end
18'd96601: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=64;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12258;
 end   
18'd96602: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=37;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd96603: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=50;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd96604: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=10;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd96605: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=91;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd96606: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd96607: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd96608: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd96609: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd96610: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd96742: begin  
rid<=1;
end
18'd96743: begin  
end
18'd96744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd96745: begin  
rid<=0;
end
18'd96801: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=3;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7139;
 end   
18'd96802: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=64;
   mapp<=21;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9702;
 end   
18'd96803: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=45;
   mapp<=18;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=11698;
 end   
18'd96804: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=49;
   mapp<=98;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=11776;
 end   
18'd96805: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=83;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=7117;
 end   
18'd96806: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=33;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=10162;
 end   
18'd96807: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=95;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=7493;
 end   
18'd96808: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd96809: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd96810: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd96811: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd96812: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd96813: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7139;
 end   
18'd96814: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7139;
 end   
18'd96942: begin  
rid<=1;
end
18'd96943: begin  
end
18'd96944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd96945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd96946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd96947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd96948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd96949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd96950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd96951: begin  
rid<=0;
end
18'd97001: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=6;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6005;
 end   
18'd97002: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=87;
   mapp<=44;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7124;
 end   
18'd97003: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=35;
   mapp<=55;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=7863;
 end   
18'd97004: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=59;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=9275;
 end   
18'd97005: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=68;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=7878;
 end   
18'd97006: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=85;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=3027;
 end   
18'd97007: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=1;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=7627;
 end   
18'd97008: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd97009: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd97010: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd97011: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd97012: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd97142: begin  
rid<=1;
end
18'd97143: begin  
end
18'd97144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd97145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd97146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd97147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd97148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd97149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd97150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd97151: begin  
rid<=0;
end
18'd97201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=25;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3889;
 end   
18'd97202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=24;
   mapp<=51;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3148;
 end   
18'd97203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=46;
   mapp<=40;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=3058;
 end   
18'd97204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=3208;
 end   
18'd97205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=38;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=3715;
 end   
18'd97206: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=31;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd97207: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=21;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd97208: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd97209: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd97210: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd97342: begin  
rid<=1;
end
18'd97343: begin  
end
18'd97344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd97345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd97346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd97347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd97348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd97349: begin  
rid<=0;
end
18'd97401: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=67;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=17413;
 end   
18'd97402: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=19;
   mapp<=15;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10079;
 end   
18'd97403: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=74;
   mapp<=44;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=14585;
 end   
18'd97404: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=87;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd97405: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=30;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd97406: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=45;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd97407: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd97408: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=44;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd97409: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd97410: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd97411: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd97412: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd97413: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17413;
 end   
18'd97414: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17413;
 end   
18'd97542: begin  
rid<=1;
end
18'd97543: begin  
end
18'd97544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd97545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd97546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd97547: begin  
rid<=0;
end
18'd97601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=11;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5655;
 end   
18'd97602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=29;
   mapp<=15;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8328;
 end   
18'd97603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=24;
   mapp<=21;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9733;
 end   
18'd97604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=59;
   mapp<=2;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=11763;
 end   
18'd97605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=83;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd97606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=65;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd97607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd97608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd97609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd97610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd97611: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd97612: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd97613: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5655;
 end   
18'd97614: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5655;
 end   
18'd97615: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5655;
 end   
18'd97742: begin  
rid<=1;
end
18'd97743: begin  
end
18'd97744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd97745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd97746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd97747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd97748: begin  
rid<=0;
end
18'd97801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=90;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10566;
 end   
18'd97802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=84;
   mapp<=91;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=16426;
 end   
18'd97803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=6;
   mapp<=97;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=10268;
 end   
18'd97804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=13;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=7680;
 end   
18'd97805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=71;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=14026;
 end   
18'd97806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd97807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd97808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd97809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd97810: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd97942: begin  
rid<=1;
end
18'd97943: begin  
end
18'd97944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd97945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd97946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd97947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd97948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd97949: begin  
rid<=0;
end
18'd98001: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=79;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15487;
 end   
18'd98002: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=98;
   mapp<=66;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10542;
 end   
18'd98003: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=67;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd98004: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=45;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd98005: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=3;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd98006: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=30;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd98007: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=20;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd98008: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=25;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd98009: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd98010: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd98011: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd98012: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd98013: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15487;
 end   
18'd98014: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15487;
 end   
18'd98015: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15487;
 end   
18'd98142: begin  
rid<=1;
end
18'd98143: begin  
end
18'd98144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd98145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd98146: begin  
rid<=0;
end
18'd98201: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=24;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5578;
 end   
18'd98202: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=92;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10528;
 end   
18'd98203: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=18;
   mapp<=87;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=11150;
 end   
18'd98204: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=93;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=5610;
 end   
18'd98205: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd98206: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd98207: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd98208: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd98209: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd98342: begin  
rid<=1;
end
18'd98343: begin  
end
18'd98344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd98345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd98346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd98347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd98348: begin  
rid<=0;
end
18'd98401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=19;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=26027;
 end   
18'd98402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=7;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd98403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=71;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd98404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=22;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd98405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=61;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd98406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=91;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd98407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=52;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd98408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=51;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd98409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd98410: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd98411: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd98412: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd98413: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26027;
 end   
18'd98414: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26027;
 end   
18'd98415: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26027;
 end   
18'd98416: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26027;
 end   
18'd98542: begin  
rid<=1;
end
18'd98543: begin  
end
18'd98544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd98545: begin  
rid<=0;
end
18'd98601: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=28;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7601;
 end   
18'd98602: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=35;
   mapp<=80;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7830;
 end   
18'd98603: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=53;
   mapp<=61;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5222;
 end   
18'd98604: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=65;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=2655;
 end   
18'd98605: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd98606: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd98607: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd98608: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd98609: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd98742: begin  
rid<=1;
end
18'd98743: begin  
end
18'd98744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd98745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd98746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd98747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd98748: begin  
rid<=0;
end
18'd98801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=61;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=18197;
 end   
18'd98802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=42;
   mapp<=57;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=20151;
 end   
18'd98803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=31;
   mapp<=89;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=18732;
 end   
18'd98804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=60;
   mapp<=92;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=20732;
 end   
18'd98805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=99;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=17825;
 end   
18'd98806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=38;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd98807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=80;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd98808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=20;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd98809: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=45;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd98810: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=29;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd98811: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd98812: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd98813: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18197;
 end   
18'd98814: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18197;
 end   
18'd98815: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18197;
 end   
18'd98816: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18197;
 end   
18'd98942: begin  
rid<=1;
end
18'd98943: begin  
end
18'd98944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd98945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd98946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd98947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd98948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd98949: begin  
rid<=0;
end
18'd99001: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=64;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=18219;
 end   
18'd99002: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=41;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd99003: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=99;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd99004: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=36;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd99005: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=65;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd99006: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=33;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd99007: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=29;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd99008: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd99009: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd99010: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd99011: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd99012: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd99013: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18219;
 end   
18'd99014: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18219;
 end   
18'd99142: begin  
rid<=1;
end
18'd99143: begin  
end
18'd99144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd99145: begin  
rid<=0;
end
18'd99201: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=6;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=20166;
 end   
18'd99202: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=10;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd99203: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=63;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd99204: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=48;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd99205: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=90;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd99206: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=69;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd99207: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=44;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd99208: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=99;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd99209: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd99210: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd99211: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd99212: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd99213: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20166;
 end   
18'd99214: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20166;
 end   
18'd99215: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20166;
 end   
18'd99216: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20166;
 end   
18'd99342: begin  
rid<=1;
end
18'd99343: begin  
end
18'd99344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd99345: begin  
rid<=0;
end
18'd99401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=6;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1603;
 end   
18'd99402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=11;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd99403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=14;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd99404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd99405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd99406: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd99542: begin  
rid<=1;
end
18'd99543: begin  
end
18'd99544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd99545: begin  
rid<=0;
end
18'd99601: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=34;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15704;
 end   
18'd99602: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=76;
   mapp<=87;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=15107;
 end   
18'd99603: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=15;
   mapp<=80;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=15808;
 end   
18'd99604: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=18;
   mapp<=85;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=18708;
 end   
18'd99605: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=84;
   mapp<=64;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=17920;
 end   
18'd99606: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=47;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd99607: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=48;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd99608: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=47;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd99609: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=55;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd99610: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd99611: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd99612: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd99613: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15704;
 end   
18'd99614: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15704;
 end   
18'd99742: begin  
rid<=1;
end
18'd99743: begin  
end
18'd99744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd99745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd99746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd99747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd99748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd99749: begin  
rid<=0;
end
18'd99801: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=4;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14992;
 end   
18'd99802: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=29;
   mapp<=27;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=12855;
 end   
18'd99803: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=15;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd99804: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=65;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd99805: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=50;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd99806: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=32;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd99807: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=83;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd99808: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=19;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd99809: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd99810: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd99811: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd99812: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd99813: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14992;
 end   
18'd99814: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14992;
 end   
18'd99815: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14992;
 end   
18'd99816: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14992;
 end   
18'd99817: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14992;
 end   
18'd99942: begin  
rid<=1;
end
18'd99943: begin  
end
18'd99944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd99945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd99946: begin  
rid<=0;
end
18'd100001: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=6;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4245;
 end   
18'd100002: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=20;
   mapp<=38;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6254;
 end   
18'd100003: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=70;
   mapp<=41;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=7619;
 end   
18'd100004: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=49;
   mapp<=3;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=5260;
 end   
18'd100005: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=5;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=4801;
 end   
18'd100006: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=24;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=8705;
 end   
18'd100007: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=78;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd100008: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=87;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd100009: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=84;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd100010: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd100011: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd100012: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd100013: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=4245;
 end   
18'd100142: begin  
rid<=1;
end
18'd100143: begin  
end
18'd100144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd100145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd100146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd100147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd100148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd100149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd100150: begin  
rid<=0;
end
18'd100201: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=38;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4819;
 end   
18'd100202: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=15;
   mapp<=73;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1626;
 end   
18'd100203: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=2;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=3209;
 end   
18'd100204: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=41;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=10253;
 end   
18'd100205: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=85;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=12969;
 end   
18'd100206: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=63;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=7027;
 end   
18'd100207: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=11;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=5956;
 end   
18'd100208: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=66;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd100209: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd100210: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd100342: begin  
rid<=1;
end
18'd100343: begin  
end
18'd100344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd100345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd100346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd100347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd100348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd100349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd100350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd100351: begin  
rid<=0;
end
18'd100401: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=12;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4164;
 end   
18'd100402: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=56;
   mapp<=65;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5546;
 end   
18'd100403: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=2;
   mapp<=82;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5658;
 end   
18'd100404: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=82;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=2820;
 end   
18'd100405: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=31;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=2552;
 end   
18'd100406: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd100407: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd100408: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd100409: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd100410: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd100542: begin  
rid<=1;
end
18'd100543: begin  
end
18'd100544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd100545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd100546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd100547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd100548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd100549: begin  
rid<=0;
end
18'd100601: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=38;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3316;
 end   
18'd100602: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=24;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5232;
 end   
18'd100603: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=64;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=2812;
 end   
18'd100604: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=15;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=2832;
 end   
18'd100605: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=93;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=3742;
 end   
18'd100606: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=7;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=1204;
 end   
18'd100607: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=37;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=1898;
 end   
18'd100608: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd100609: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd100610: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd100742: begin  
rid<=1;
end
18'd100743: begin  
end
18'd100744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd100745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd100746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd100747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd100748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd100749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd100750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd100751: begin  
rid<=0;
end
18'd100801: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=37;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9888;
 end   
18'd100802: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=60;
   mapp<=28;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=12433;
 end   
18'd100803: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=49;
   mapp<=59;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9168;
 end   
18'd100804: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=23;
   mapp<=83;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=7858;
 end   
18'd100805: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=83;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd100806: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=5;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd100807: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=47;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd100808: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=13;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd100809: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd100810: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd100811: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd100812: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd100813: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9888;
 end   
18'd100942: begin  
rid<=1;
end
18'd100943: begin  
end
18'd100944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd100945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd100946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd100947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd100948: begin  
rid<=0;
end
18'd101001: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=39;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2289;
 end   
18'd101002: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=57;
   mapp<=34;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1336;
 end   
18'd101003: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=4010;
 end   
18'd101004: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd101005: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd101006: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd101142: begin  
rid<=1;
end
18'd101143: begin  
end
18'd101144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd101145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd101146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd101147: begin  
rid<=0;
end
18'd101201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=35;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14472;
 end   
18'd101202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=83;
   mapp<=92;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13740;
 end   
18'd101203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=27;
   mapp<=22;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=15735;
 end   
18'd101204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=99;
   mapp<=33;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=17192;
 end   
18'd101205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=61;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd101206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=90;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd101207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=35;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd101208: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd101209: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd101210: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd101211: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd101342: begin  
rid<=1;
end
18'd101343: begin  
end
18'd101344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd101345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd101346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd101347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd101348: begin  
rid<=0;
end
18'd101401: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=6;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=438;
 end   
18'd101402: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=85;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6215;
 end   
18'd101403: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=45;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=3305;
 end   
18'd101404: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=9;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=687;
 end   
18'd101405: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=36;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=2668;
 end   
18'd101406: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=81;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=5963;
 end   
18'd101407: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=39;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=2907;
 end   
18'd101408: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=99;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=7297;
 end   
18'd101409: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd101542: begin  
rid<=1;
end
18'd101543: begin  
end
18'd101544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd101545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd101546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd101547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd101548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd101549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd101550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd101551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd101552: begin  
rid<=0;
end
18'd101601: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=33;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4123;
 end   
18'd101602: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=52;
   mapp<=19;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5005;
 end   
18'd101603: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=84;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=4196;
 end   
18'd101604: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=27;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=3781;
 end   
18'd101605: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd101606: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd101607: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd101608: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd101609: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd101742: begin  
rid<=1;
end
18'd101743: begin  
end
18'd101744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd101745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd101746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd101747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd101748: begin  
rid<=0;
end
18'd101801: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=49;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=29700;
 end   
18'd101802: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=90;
   mapp<=75;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=32360;
 end   
18'd101803: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=46;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd101804: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=98;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd101805: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=67;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd101806: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=46;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd101807: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=9;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd101808: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=80;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd101809: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=79;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd101810: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd101811: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd101812: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd101813: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29700;
 end   
18'd101814: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29700;
 end   
18'd101815: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29700;
 end   
18'd101816: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29700;
 end   
18'd101817: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29700;
 end   
18'd101818: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29700;
 end   
18'd101819: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29700;
 end   
18'd101942: begin  
rid<=1;
end
18'd101943: begin  
end
18'd101944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd101945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd101946: begin  
rid<=0;
end
18'd102001: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=55;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8226;
 end   
18'd102002: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=32;
   mapp<=38;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9094;
 end   
18'd102003: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=65;
   mapp<=25;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=10738;
 end   
18'd102004: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=18;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd102005: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=20;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd102006: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=37;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd102007: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=64;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd102008: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=9;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd102009: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=3;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd102010: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd102011: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd102012: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd102013: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8226;
 end   
18'd102014: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8226;
 end   
18'd102015: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8226;
 end   
18'd102016: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8226;
 end   
18'd102142: begin  
rid<=1;
end
18'd102143: begin  
end
18'd102144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd102145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd102146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd102147: begin  
rid<=0;
end
18'd102201: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=24;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13614;
 end   
18'd102202: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=83;
   mapp<=1;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=12878;
 end   
18'd102203: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=98;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd102204: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=40;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd102205: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=31;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd102206: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=70;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd102207: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=54;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd102208: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=35;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd102209: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd102210: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd102211: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd102212: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd102213: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13614;
 end   
18'd102214: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13614;
 end   
18'd102215: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13614;
 end   
18'd102342: begin  
rid<=1;
end
18'd102343: begin  
end
18'd102344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd102345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd102346: begin  
rid<=0;
end
18'd102401: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=30;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1767;
 end   
18'd102402: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=18;
   mapp<=14;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2566;
 end   
18'd102403: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=32;
   mapp<=32;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=4407;
 end   
18'd102404: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=13;
   mapp<=17;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=3903;
 end   
18'd102405: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=90;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=3323;
 end   
18'd102406: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=61;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=2456;
 end   
18'd102407: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=32;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd102408: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=35;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd102409: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=17;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd102410: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd102411: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd102412: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd102413: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=1767;
 end   
18'd102542: begin  
rid<=1;
end
18'd102543: begin  
end
18'd102544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd102545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd102546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd102547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd102548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd102549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd102550: begin  
rid<=0;
end
18'd102601: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=46;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6056;
 end   
18'd102602: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=70;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4980;
 end   
18'd102603: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=88;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd102604: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=94;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd102605: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=8;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd102606: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd102607: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd102608: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd102609: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd102742: begin  
rid<=1;
end
18'd102743: begin  
end
18'd102744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd102745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd102746: begin  
rid<=0;
end
18'd102801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=5;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4135;
 end   
18'd102802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=50;
   mapp<=75;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7010;
 end   
18'd102803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=42;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd102804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd102805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd102942: begin  
rid<=1;
end
18'd102943: begin  
end
18'd102944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd102945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd102946: begin  
rid<=0;
end
18'd103001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=71;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10394;
 end   
18'd103002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=22;
   mapp<=24;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6312;
 end   
18'd103003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=44;
   mapp<=79;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9435;
 end   
18'd103004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd103005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd103006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd103007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd103008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd103142: begin  
rid<=1;
end
18'd103143: begin  
end
18'd103144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd103145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd103146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd103147: begin  
rid<=0;
end
18'd103201: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=41;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9980;
 end   
18'd103202: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=17;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13883;
 end   
18'd103203: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=68;
   mapp<=52;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=14951;
 end   
18'd103204: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=65;
   mapp<=74;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=15519;
 end   
18'd103205: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=77;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=12271;
 end   
18'd103206: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=97;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=12360;
 end   
18'd103207: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd103208: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd103209: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd103210: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd103211: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd103212: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd103213: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9980;
 end   
18'd103342: begin  
rid<=1;
end
18'd103343: begin  
end
18'd103344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd103345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd103346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd103347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd103348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd103349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd103350: begin  
rid<=0;
end
18'd103401: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=92;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=17348;
 end   
18'd103402: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=35;
   mapp<=14;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=15576;
 end   
18'd103403: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=30;
   mapp<=83;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12913;
 end   
18'd103404: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=34;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd103405: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=20;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd103406: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=28;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd103407: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=88;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd103408: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=24;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd103409: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=34;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd103410: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=33;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd103411: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=3;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd103412: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd103413: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17348;
 end   
18'd103414: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17348;
 end   
18'd103415: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17348;
 end   
18'd103416: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17348;
 end   
18'd103417: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17348;
 end   
18'd103418: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17348;
 end   
18'd103419: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17348;
 end   
18'd103420: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17348;
 end   
18'd103542: begin  
rid<=1;
end
18'd103543: begin  
end
18'd103544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd103545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd103546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd103547: begin  
rid<=0;
end
18'd103601: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=31;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16236;
 end   
18'd103602: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=65;
   mapp<=60;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=15642;
 end   
18'd103603: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=26;
   mapp<=65;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=15321;
 end   
18'd103604: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=62;
   mapp<=30;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=13846;
 end   
18'd103605: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=63;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd103606: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=78;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd103607: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=19;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd103608: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd103609: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd103610: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd103611: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd103612: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd103613: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16236;
 end   
18'd103614: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16236;
 end   
18'd103615: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16236;
 end   
18'd103616: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16236;
 end   
18'd103617: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16236;
 end   
18'd103742: begin  
rid<=1;
end
18'd103743: begin  
end
18'd103744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd103745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd103746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd103747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd103748: begin  
rid<=0;
end
18'd103801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=39;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=23316;
 end   
18'd103802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=39;
   mapp<=76;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=20291;
 end   
18'd103803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=52;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd103804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=30;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd103805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=74;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd103806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=81;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd103807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=42;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd103808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=18;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd103809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd103810: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd103811: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd103812: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd103813: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23316;
 end   
18'd103814: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23316;
 end   
18'd103815: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23316;
 end   
18'd103942: begin  
rid<=1;
end
18'd103943: begin  
end
18'd103944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd103945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd103946: begin  
rid<=0;
end
18'd104001: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=34;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1156;
 end   
18'd104002: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=6;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=214;
 end   
18'd104003: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=80;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=2740;
 end   
18'd104004: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=90;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=3090;
 end   
18'd104005: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=23;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=822;
 end   
18'd104006: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=99;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=3416;
 end   
18'd104007: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=68;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=2372;
 end   
18'd104008: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=85;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=2960;
 end   
18'd104009: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd104142: begin  
rid<=1;
end
18'd104143: begin  
end
18'd104144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd104145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd104146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd104147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd104148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd104149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd104150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd104151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd104152: begin  
rid<=0;
end
18'd104201: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=0;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=152;
 end   
18'd104202: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=19;
   mapp<=8;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=990;
 end   
18'd104203: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=18;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1204;
 end   
18'd104204: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=49;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=2562;
 end   
18'd104205: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=47;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=2748;
 end   
18'd104206: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=80;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=4362;
 end   
18'd104207: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=99;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=4800;
 end   
18'd104208: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=48;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=2854;
 end   
18'd104209: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=84;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=3928;
 end   
18'd104210: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=19;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd104211: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd104212: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd104342: begin  
rid<=1;
end
18'd104343: begin  
end
18'd104344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd104345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd104346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd104347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd104348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd104349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd104350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd104351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd104352: begin  
check<=expctdoutput[8]-outcheck;
end
18'd104353: begin  
rid<=0;
end
18'd104401: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=22;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11857;
 end   
18'd104402: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=45;
   mapp<=70;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=14319;
 end   
18'd104403: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=40;
   mapp<=97;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=14866;
 end   
18'd104404: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=27;
   mapp<=33;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=19371;
 end   
18'd104405: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=50;
   mapp<=40;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=20006;
 end   
18'd104406: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=82;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=23009;
 end   
18'd104407: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=47;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd104408: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=99;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd104409: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=50;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd104410: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=30;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd104411: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd104412: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd104413: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11857;
 end   
18'd104414: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11857;
 end   
18'd104415: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11857;
 end   
18'd104542: begin  
rid<=1;
end
18'd104543: begin  
end
18'd104544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd104545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd104546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd104547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd104548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd104549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd104550: begin  
rid<=0;
end
18'd104601: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=39;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1544;
 end   
18'd104602: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=67;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3622;
 end   
18'd104603: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=51;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=7503;
 end   
18'd104604: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd104605: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd104606: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd104742: begin  
rid<=1;
end
18'd104743: begin  
end
18'd104744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd104745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd104746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd104747: begin  
rid<=0;
end
18'd104801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=66;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=18203;
 end   
18'd104802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=33;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=21009;
 end   
18'd104803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=43;
   mapp<=73;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=15720;
 end   
18'd104804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=72;
   mapp<=16;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=19555;
 end   
18'd104805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=14;
   mapp<=57;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=16156;
 end   
18'd104806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=98;
   mapp<=86;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=14150;
 end   
18'd104807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=71;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd104808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd104809: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=61;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd104810: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=9;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd104811: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=20;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd104812: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd104813: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18203;
 end   
18'd104814: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18203;
 end   
18'd104815: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18203;
 end   
18'd104816: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18203;
 end   
18'd104817: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18203;
 end   
18'd104942: begin  
rid<=1;
end
18'd104943: begin  
end
18'd104944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd104945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd104946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd104947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd104948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd104949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd104950: begin  
rid<=0;
end
18'd105001: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=28;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8202;
 end   
18'd105002: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=91;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd105003: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=97;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd105004: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd105005: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd105006: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd105142: begin  
rid<=1;
end
18'd105143: begin  
end
18'd105144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd105145: begin  
rid<=0;
end
18'd105201: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=90;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2070;
 end   
18'd105202: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=10;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=910;
 end   
18'd105203: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=71;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=6410;
 end   
18'd105204: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=78;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=7050;
 end   
18'd105205: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=93;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=8410;
 end   
18'd105206: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd105342: begin  
rid<=1;
end
18'd105343: begin  
end
18'd105344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd105345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd105346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd105347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd105348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd105349: begin  
rid<=0;
end
18'd105401: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=88;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11996;
 end   
18'd105402: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=22;
   mapp<=47;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13123;
 end   
18'd105403: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=77;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd105404: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=19;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd105405: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=83;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd105406: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd105407: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd105408: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd105409: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd105410: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd105411: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd105542: begin  
rid<=1;
end
18'd105543: begin  
end
18'd105544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd105545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd105546: begin  
rid<=0;
end
18'd105601: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=97;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=23822;
 end   
18'd105602: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=66;
   mapp<=46;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=23769;
 end   
18'd105603: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=60;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd105604: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=91;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd105605: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=73;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd105606: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd105607: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd105608: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd105609: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd105610: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd105611: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd105742: begin  
rid<=1;
end
18'd105743: begin  
end
18'd105744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd105745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd105746: begin  
rid<=0;
end
18'd105801: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=38;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=228;
 end   
18'd105802: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=96;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=586;
 end   
18'd105803: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=18;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=128;
 end   
18'd105804: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=62;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=402;
 end   
18'd105805: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=44;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=304;
 end   
18'd105806: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=26;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=206;
 end   
18'd105807: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=15;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=150;
 end   
18'd105808: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=93;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=628;
 end   
18'd105809: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd105942: begin  
rid<=1;
end
18'd105943: begin  
end
18'd105944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd105945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd105946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd105947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd105948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd105949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd105950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd105951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd105952: begin  
rid<=0;
end
18'd106001: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=29;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16870;
 end   
18'd106002: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=94;
   mapp<=18;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=18897;
 end   
18'd106003: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=37;
   mapp<=69;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=18849;
 end   
18'd106004: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=95;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd106005: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=30;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd106006: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=49;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd106007: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd106008: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd106009: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd106010: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd106011: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd106012: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd106013: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16870;
 end   
18'd106014: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16870;
 end   
18'd106142: begin  
rid<=1;
end
18'd106143: begin  
end
18'd106144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd106145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd106146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd106147: begin  
rid<=0;
end
18'd106201: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=55;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=18675;
 end   
18'd106202: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=61;
   mapp<=61;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=15007;
 end   
18'd106203: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=51;
   mapp<=3;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=14285;
 end   
18'd106204: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=10;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd106205: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=77;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd106206: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=76;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd106207: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=39;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd106208: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=22;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd106209: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd106210: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd106211: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd106212: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd106213: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18675;
 end   
18'd106214: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18675;
 end   
18'd106215: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18675;
 end   
18'd106216: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18675;
 end   
18'd106217: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18675;
 end   
18'd106218: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18675;
 end   
18'd106342: begin  
rid<=1;
end
18'd106343: begin  
end
18'd106344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd106345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd106346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd106347: begin  
rid<=0;
end
18'd106401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=12;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2601;
 end   
18'd106402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=23;
   mapp<=49;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4537;
 end   
18'd106403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=14;
   mapp<=23;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5027;
 end   
18'd106404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=71;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=7698;
 end   
18'd106405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=8;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd106406: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=20;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd106407: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd106408: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd106409: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd106542: begin  
rid<=1;
end
18'd106543: begin  
end
18'd106544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd106545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd106546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd106547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd106548: begin  
rid<=0;
end
18'd106601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=92;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9016;
 end   
18'd106602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=49;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=4518;
 end   
18'd106603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=45;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=4160;
 end   
18'd106604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=97;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=8954;
 end   
18'd106605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=66;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=6112;
 end   
18'd106606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=43;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=4006;
 end   
18'd106607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=48;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=4476;
 end   
18'd106608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd106742: begin  
rid<=1;
end
18'd106743: begin  
end
18'd106744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd106745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd106746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd106747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd106748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd106749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd106750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd106751: begin  
rid<=0;
end
18'd106801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=50;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9356;
 end   
18'd106802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=49;
   mapp<=94;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9459;
 end   
18'd106803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=51;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12479;
 end   
18'd106804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=81;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=16937;
 end   
18'd106805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=98;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=13580;
 end   
18'd106806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=45;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=11375;
 end   
18'd106807: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=75;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=11415;
 end   
18'd106808: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=45;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd106809: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd106810: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd106942: begin  
rid<=1;
end
18'd106943: begin  
end
18'd106944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd106945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd106946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd106947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd106948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd106949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd106950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd106951: begin  
rid<=0;
end
18'd107001: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=9;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15739;
 end   
18'd107002: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=41;
   mapp<=99;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=19218;
 end   
18'd107003: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=31;
   mapp<=67;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=23565;
 end   
18'd107004: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=99;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd107005: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=98;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd107006: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=74;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd107007: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd107008: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd107009: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd107010: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd107142: begin  
rid<=1;
end
18'd107143: begin  
end
18'd107144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd107145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd107146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd107147: begin  
rid<=0;
end
18'd107201: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=45;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2790;
 end   
18'd107202: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd107342: begin  
rid<=1;
end
18'd107343: begin  
end
18'd107344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd107345: begin  
rid<=0;
end
18'd107401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=17;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=29788;
 end   
18'd107402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=11;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=29758;
 end   
18'd107403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=68;
   mapp<=66;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=28571;
 end   
18'd107404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=48;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd107405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=81;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd107406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=33;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd107407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=74;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd107408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=88;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd107409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=84;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd107410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd107411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd107412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd107413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29788;
 end   
18'd107414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29788;
 end   
18'd107415: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29788;
 end   
18'd107416: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29788;
 end   
18'd107417: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29788;
 end   
18'd107418: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29788;
 end   
18'd107419: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29788;
 end   
18'd107420: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29788;
 end   
18'd107542: begin  
rid<=1;
end
18'd107543: begin  
end
18'd107544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd107545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd107546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd107547: begin  
rid<=0;
end
18'd107601: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=44;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1184;
 end   
18'd107602: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=21;
   mapp<=4;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=775;
 end   
18'd107603: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=60;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1564;
 end   
18'd107604: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=11;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=393;
 end   
18'd107605: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=22;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=794;
 end   
18'd107606: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=51;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=1325;
 end   
18'd107607: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=228;
 end   
18'd107608: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=42;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd107609: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd107610: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd107742: begin  
rid<=1;
end
18'd107743: begin  
end
18'd107744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd107745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd107746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd107747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd107748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd107749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd107750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd107751: begin  
rid<=0;
end
18'd107801: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=27;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13026;
 end   
18'd107802: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=80;
   mapp<=51;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6755;
 end   
18'd107803: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=5;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd107804: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=82;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd107805: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=25;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd107806: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd107807: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd107808: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd107809: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd107942: begin  
rid<=1;
end
18'd107943: begin  
end
18'd107944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd107945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd107946: begin  
rid<=0;
end
18'd108001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=26;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8331;
 end   
18'd108002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=86;
   mapp<=92;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4506;
 end   
18'd108003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=35;
   mapp<=9;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=3697;
 end   
18'd108004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=38;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=3758;
 end   
18'd108005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=5;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=8156;
 end   
18'd108006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=66;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=9927;
 end   
18'd108007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=66;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=10682;
 end   
18'd108008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=71;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=11036;
 end   
18'd108009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=80;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=9099;
 end   
18'd108010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd108011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd108012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd108013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8331;
 end   
18'd108014: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8331;
 end   
18'd108142: begin  
rid<=1;
end
18'd108143: begin  
end
18'd108144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd108145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd108146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd108147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd108148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd108149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd108150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd108151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd108152: begin  
check<=expctdoutput[8]-outcheck;
end
18'd108153: begin  
rid<=0;
end
18'd108201: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=7;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14290;
 end   
18'd108202: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=87;
   mapp<=76;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11484;
 end   
18'd108203: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=27;
   mapp<=92;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9329;
 end   
18'd108204: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=20;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd108205: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=5;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd108206: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=27;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd108207: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=37;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd108208: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=10;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd108209: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=83;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd108210: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd108211: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd108212: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd108213: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14290;
 end   
18'd108214: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14290;
 end   
18'd108215: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14290;
 end   
18'd108216: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14290;
 end   
18'd108342: begin  
rid<=1;
end
18'd108343: begin  
end
18'd108344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd108345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd108346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd108347: begin  
rid<=0;
end
18'd108401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=21;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4900;
 end   
18'd108402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=77;
   mapp<=41;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3566;
 end   
18'd108403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd108404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd108405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd108542: begin  
rid<=1;
end
18'd108543: begin  
end
18'd108544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd108545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd108546: begin  
rid<=0;
end
18'd108601: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=30;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4522;
 end   
18'd108602: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=8;
   mapp<=11;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3700;
 end   
18'd108603: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=30;
   mapp<=29;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=4669;
 end   
18'd108604: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=48;
   mapp<=53;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=6913;
 end   
18'd108605: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=32;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd108606: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=41;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd108607: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd108608: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd108609: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd108610: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd108611: begin  
  clrr<=0;
  maplen<=4;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd108742: begin  
rid<=1;
end
18'd108743: begin  
end
18'd108744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd108745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd108746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd108747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd108748: begin  
rid<=0;
end
18'd108801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=85;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16610;
 end   
18'd108802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=8;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd108803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=60;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd108804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=48;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd108805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=85;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd108806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=78;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd108807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd108808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd108809: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd108810: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd108811: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd108812: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd108942: begin  
rid<=1;
end
18'd108943: begin  
end
18'd108944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd108945: begin  
rid<=0;
end
18'd109001: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=87;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9808;
 end   
18'd109002: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=70;
   mapp<=1;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10262;
 end   
18'd109003: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=25;
   mapp<=96;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5507;
 end   
18'd109004: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=84;
   mapp<=72;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=8760;
 end   
18'd109005: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=2;
   mapp<=9;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=14304;
 end   
18'd109006: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=27;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd109007: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=46;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd109008: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd109009: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=52;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd109010: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=97;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd109011: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd109012: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd109013: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9808;
 end   
18'd109014: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9808;
 end   
18'd109015: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9808;
 end   
18'd109016: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9808;
 end   
18'd109142: begin  
rid<=1;
end
18'd109143: begin  
end
18'd109144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd109145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd109146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd109147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd109148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd109149: begin  
rid<=0;
end
18'd109201: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=18;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5487;
 end   
18'd109202: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=73;
   mapp<=51;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10071;
 end   
18'd109203: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=57;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6575;
 end   
18'd109204: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=19;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=5615;
 end   
18'd109205: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=73;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=7959;
 end   
18'd109206: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=15;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=4988;
 end   
18'd109207: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=68;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=10957;
 end   
18'd109208: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=83;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=8714;
 end   
18'd109209: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=10;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=4069;
 end   
18'd109210: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=59;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd109211: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd109212: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd109342: begin  
rid<=1;
end
18'd109343: begin  
end
18'd109344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd109345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd109346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd109347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd109348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd109349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd109350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd109351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd109352: begin  
check<=expctdoutput[8]-outcheck;
end
18'd109353: begin  
rid<=0;
end
18'd109401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=59;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4893;
 end   
18'd109402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=18;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6981;
 end   
18'd109403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=61;
   mapp<=18;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8014;
 end   
18'd109404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=67;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=4080;
 end   
18'd109405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=3;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=6319;
 end   
18'd109406: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=66;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=6246;
 end   
18'd109407: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=38;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=5374;
 end   
18'd109408: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=26;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd109409: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=93;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd109410: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd109411: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd109412: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd109542: begin  
rid<=1;
end
18'd109543: begin  
end
18'd109544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd109545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd109546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd109547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd109548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd109549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd109550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd109551: begin  
rid<=0;
end
18'd109601: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=21;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9620;
 end   
18'd109602: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=73;
   mapp<=38;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=12809;
 end   
18'd109603: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=98;
   mapp<=57;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12349;
 end   
18'd109604: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=80;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=13296;
 end   
18'd109605: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=54;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=12846;
 end   
18'd109606: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=78;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=12805;
 end   
18'd109607: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd109608: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd109609: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd109610: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd109611: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd109742: begin  
rid<=1;
end
18'd109743: begin  
end
18'd109744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd109745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd109746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd109747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd109748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd109749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd109750: begin  
rid<=0;
end
18'd109801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=39;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7163;
 end   
18'd109802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=25;
   mapp<=45;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9816;
 end   
18'd109803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=25;
   mapp<=1;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=7610;
 end   
18'd109804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=32;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd109805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=78;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd109806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=21;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd109807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd109808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd109809: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd109810: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd109811: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd109812: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd109813: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7163;
 end   
18'd109814: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7163;
 end   
18'd109942: begin  
rid<=1;
end
18'd109943: begin  
end
18'd109944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd109945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd109946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd109947: begin  
rid<=0;
end
18'd110001: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=90;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6735;
 end   
18'd110002: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=99;
   mapp<=30;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5877;
 end   
18'd110003: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=69;
   mapp<=5;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=3117;
 end   
18'd110004: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=7;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd110005: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=53;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd110006: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd110007: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd110008: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd110142: begin  
rid<=1;
end
18'd110143: begin  
end
18'd110144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd110145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd110146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd110147: begin  
rid<=0;
end
18'd110201: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=71;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16099;
 end   
18'd110202: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=64;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=18182;
 end   
18'd110203: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=99;
   mapp<=48;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=19181;
 end   
18'd110204: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=93;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=19107;
 end   
18'd110205: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=99;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=11631;
 end   
18'd110206: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=62;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=11370;
 end   
18'd110207: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=6;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=8175;
 end   
18'd110208: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=66;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=8877;
 end   
18'd110209: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd110210: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd110211: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd110212: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd110213: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16099;
 end   
18'd110342: begin  
rid<=1;
end
18'd110343: begin  
end
18'd110344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd110345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd110346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd110347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd110348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd110349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd110350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd110351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd110352: begin  
rid<=0;
end
18'd110401: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=22;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1790;
 end   
18'd110402: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=27;
   mapp<=14;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1286;
 end   
18'd110403: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=92;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd110404: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd110405: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd110406: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd110407: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd110542: begin  
rid<=1;
end
18'd110543: begin  
end
18'd110544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd110545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd110546: begin  
rid<=0;
end
18'd110601: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=52;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16463;
 end   
18'd110602: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=17;
   mapp<=71;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=19504;
 end   
18'd110603: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=24;
   mapp<=86;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=24806;
 end   
18'd110604: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=88;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd110605: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=93;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd110606: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd110607: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd110608: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd110609: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd110610: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd110742: begin  
rid<=1;
end
18'd110743: begin  
end
18'd110744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd110745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd110746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd110747: begin  
rid<=0;
end
18'd110801: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=37;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=22437;
 end   
18'd110802: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=43;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=17916;
 end   
18'd110803: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=7;
   mapp<=46;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=18838;
 end   
18'd110804: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=70;
   mapp<=58;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=17670;
 end   
18'd110805: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=49;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd110806: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=46;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd110807: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=39;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd110808: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=52;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd110809: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd110810: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd110811: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd110812: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd110813: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22437;
 end   
18'd110814: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22437;
 end   
18'd110815: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22437;
 end   
18'd110816: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22437;
 end   
18'd110817: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22437;
 end   
18'd110818: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22437;
 end   
18'd110819: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22437;
 end   
18'd110942: begin  
rid<=1;
end
18'd110943: begin  
end
18'd110944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd110945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd110946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd110947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd110948: begin  
rid<=0;
end
18'd111001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=99;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15884;
 end   
18'd111002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=16;
   mapp<=76;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=16391;
 end   
18'd111003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=74;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd111004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=56;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd111005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=77;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd111006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=72;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd111007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd111008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd111009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd111010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd111011: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd111142: begin  
rid<=1;
end
18'd111143: begin  
end
18'd111144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd111145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd111146: begin  
rid<=0;
end
18'd111201: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=32;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3594;
 end   
18'd111202: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=58;
   mapp<=9;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6370;
 end   
18'd111203: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=88;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8864;
 end   
18'd111204: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=44;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=4290;
 end   
18'd111205: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=4;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=694;
 end   
18'd111206: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=30;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=3173;
 end   
18'd111207: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=27;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=3093;
 end   
18'd111208: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=49;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd111209: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd111210: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd111342: begin  
rid<=1;
end
18'd111343: begin  
end
18'd111344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd111345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd111346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd111347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd111348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd111349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd111350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd111351: begin  
rid<=0;
end
18'd111401: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=62;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14064;
 end   
18'd111402: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=80;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd111403: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=18;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd111404: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=28;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd111405: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=89;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd111406: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=13;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd111407: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=41;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd111408: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd111409: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd111410: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd111411: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd111412: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd111413: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14064;
 end   
18'd111414: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14064;
 end   
18'd111542: begin  
rid<=1;
end
18'd111543: begin  
end
18'd111544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd111545: begin  
rid<=0;
end
18'd111601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=52;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3923;
 end   
18'd111602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=57;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3892;
 end   
18'd111603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=1;
   mapp<=31;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=3659;
 end   
18'd111604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=35;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=3756;
 end   
18'd111605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=32;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=6460;
 end   
18'd111606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=82;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=9038;
 end   
18'd111607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=82;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=7218;
 end   
18'd111608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd111609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd111610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd111611: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd111612: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd111742: begin  
rid<=1;
end
18'd111743: begin  
end
18'd111744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd111745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd111746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd111747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd111748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd111749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd111750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd111751: begin  
rid<=0;
end
18'd111801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=82;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7114;
 end   
18'd111802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=12;
   mapp<=94;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7946;
 end   
18'd111803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=19;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=1890;
 end   
18'd111804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=26;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=3158;
 end   
18'd111805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=83;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=7242;
 end   
18'd111806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd111807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd111808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd111942: begin  
rid<=1;
end
18'd111943: begin  
end
18'd111944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd111945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd111946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd111947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd111948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd111949: begin  
rid<=0;
end
18'd112001: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=24;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1788;
 end   
18'd112002: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=45;
   mapp<=12;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3502;
 end   
18'd112003: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=96;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5036;
 end   
18'd112004: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=2;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=1010;
 end   
18'd112005: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=73;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=4532;
 end   
18'd112006: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=58;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=3126;
 end   
18'd112007: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=5;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd112008: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd112009: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd112142: begin  
rid<=1;
end
18'd112143: begin  
end
18'd112144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd112145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd112146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd112147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd112148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd112149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd112150: begin  
rid<=0;
end
18'd112201: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=50;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6220;
 end   
18'd112202: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=70;
   mapp<=81;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7260;
 end   
18'd112203: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=80;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5193;
 end   
18'd112204: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=53;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=2800;
 end   
18'd112205: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=27;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=5116;
 end   
18'd112206: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=59;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=1995;
 end   
18'd112207: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=16;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=8093;
 end   
18'd112208: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=97;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd112209: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd112210: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd112342: begin  
rid<=1;
end
18'd112343: begin  
end
18'd112344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd112345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd112346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd112347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd112348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd112349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd112350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd112351: begin  
rid<=0;
end
18'd112401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=52;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9672;
 end   
18'd112402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=13;
   mapp<=81;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11702;
 end   
18'd112403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=71;
   mapp<=65;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=17233;
 end   
18'd112404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=76;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=17658;
 end   
18'd112405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=86;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=15386;
 end   
18'd112406: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=74;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=11815;
 end   
18'd112407: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=42;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=7200;
 end   
18'd112408: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=41;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd112409: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=9;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd112410: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd112411: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd112412: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd112542: begin  
rid<=1;
end
18'd112543: begin  
end
18'd112544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd112545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd112546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd112547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd112548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd112549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd112550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd112551: begin  
rid<=0;
end
18'd112601: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=48;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6168;
 end   
18'd112602: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=92;
   mapp<=42;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5938;
 end   
18'd112603: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=36;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=2588;
 end   
18'd112604: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=20;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd112605: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd112606: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd112742: begin  
rid<=1;
end
18'd112743: begin  
end
18'd112744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd112745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd112746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd112747: begin  
rid<=0;
end
18'd112801: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=5;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=20269;
 end   
18'd112802: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=81;
   mapp<=81;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=22048;
 end   
18'd112803: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=68;
   mapp<=38;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=19526;
 end   
18'd112804: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=14;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd112805: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=1;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd112806: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=16;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd112807: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=94;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd112808: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=67;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd112809: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=45;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd112810: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=67;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd112811: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=39;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd112812: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd112813: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20269;
 end   
18'd112814: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20269;
 end   
18'd112815: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20269;
 end   
18'd112816: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20269;
 end   
18'd112817: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20269;
 end   
18'd112818: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20269;
 end   
18'd112819: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20269;
 end   
18'd112820: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20269;
 end   
18'd112942: begin  
rid<=1;
end
18'd112943: begin  
end
18'd112944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd112945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd112946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd112947: begin  
rid<=0;
end
18'd113001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=17;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15235;
 end   
18'd113002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=24;
   mapp<=44;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=18866;
 end   
18'd113003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=49;
   mapp<=99;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=22981;
 end   
18'd113004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=86;
   mapp<=25;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=18618;
 end   
18'd113005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=74;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd113006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=57;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd113007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=85;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd113008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=15;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd113009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd113010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd113011: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd113012: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd113013: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15235;
 end   
18'd113142: begin  
rid<=1;
end
18'd113143: begin  
end
18'd113144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd113145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd113146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd113147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd113148: begin  
rid<=0;
end
18'd113201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=70;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9221;
 end   
18'd113202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=62;
   mapp<=82;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11897;
 end   
18'd113203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=91;
   mapp<=11;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6161;
 end   
18'd113204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=28;
   mapp<=37;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=9556;
 end   
18'd113205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=61;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=6722;
 end   
18'd113206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=12;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=9118;
 end   
18'd113207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=96;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=11318;
 end   
18'd113208: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=76;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=5615;
 end   
18'd113209: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd113210: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=58;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd113211: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=71;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd113212: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd113213: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9221;
 end   
18'd113214: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9221;
 end   
18'd113215: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9221;
 end   
18'd113342: begin  
rid<=1;
end
18'd113343: begin  
end
18'd113344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd113345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd113346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd113347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd113348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd113349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd113350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd113351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd113352: begin  
rid<=0;
end
18'd113401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=58;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6270;
 end   
18'd113402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=28;
   mapp<=98;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7136;
 end   
18'd113403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=45;
   mapp<=50;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=7026;
 end   
18'd113404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=42;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=7678;
 end   
18'd113405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd113406: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=60;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd113407: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd113408: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd113409: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd113542: begin  
rid<=1;
end
18'd113543: begin  
end
18'd113544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd113545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd113546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd113547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd113548: begin  
rid<=0;
end
18'd113601: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=95;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8835;
 end   
18'd113602: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=4;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=382;
 end   
18'd113603: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=13;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1229;
 end   
18'd113604: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd113742: begin  
rid<=1;
end
18'd113743: begin  
end
18'd113744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd113745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd113746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd113747: begin  
rid<=0;
end
18'd113801: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=95;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=380;
 end   
18'd113802: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=21;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=94;
 end   
18'd113803: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=48;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=212;
 end   
18'd113804: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=68;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=302;
 end   
18'd113805: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd113942: begin  
rid<=1;
end
18'd113943: begin  
end
18'd113944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd113945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd113946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd113947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd113948: begin  
rid<=0;
end
18'd114001: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=32;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3634;
 end   
18'd114002: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=19;
   mapp<=38;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3145;
 end   
18'd114003: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=37;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5895;
 end   
18'd114004: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=66;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=7252;
 end   
18'd114005: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=32;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=5308;
 end   
18'd114006: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=62;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=6984;
 end   
18'd114007: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd114008: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd114009: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd114142: begin  
rid<=1;
end
18'd114143: begin  
end
18'd114144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd114145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd114146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd114147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd114148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd114149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd114150: begin  
rid<=0;
end
18'd114201: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=6;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6231;
 end   
18'd114202: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=11;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7174;
 end   
18'd114203: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=97;
   mapp<=11;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9581;
 end   
18'd114204: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=37;
   mapp<=14;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=9957;
 end   
18'd114205: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=2;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd114206: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=15;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd114207: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=63;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd114208: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=17;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd114209: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd114210: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd114211: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd114212: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd114213: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6231;
 end   
18'd114214: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6231;
 end   
18'd114215: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6231;
 end   
18'd114216: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6231;
 end   
18'd114217: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6231;
 end   
18'd114218: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6231;
 end   
18'd114219: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6231;
 end   
18'd114342: begin  
rid<=1;
end
18'd114343: begin  
end
18'd114344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd114345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd114346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd114347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd114348: begin  
rid<=0;
end
18'd114401: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=87;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9211;
 end   
18'd114402: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=12;
   mapp<=43;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9004;
 end   
18'd114403: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=12;
   mapp<=38;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=13966;
 end   
18'd114404: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=22;
   mapp<=82;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=13449;
 end   
18'd114405: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=37;
   mapp<=54;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=10195;
 end   
18'd114406: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=74;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=12271;
 end   
18'd114407: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=91;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd114408: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=8;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd114409: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=18;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd114410: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=51;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd114411: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd114412: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd114413: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9211;
 end   
18'd114414: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9211;
 end   
18'd114415: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9211;
 end   
18'd114542: begin  
rid<=1;
end
18'd114543: begin  
end
18'd114544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd114545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd114546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd114547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd114548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd114549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd114550: begin  
rid<=0;
end
18'd114601: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=29;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=18394;
 end   
18'd114602: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=21;
   mapp<=11;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10101;
 end   
18'd114603: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=87;
   mapp<=30;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=20268;
 end   
18'd114604: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=63;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd114605: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=27;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd114606: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=88;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd114607: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=77;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd114608: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=14;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd114609: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=46;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd114610: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=75;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd114611: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd114612: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd114613: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18394;
 end   
18'd114614: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18394;
 end   
18'd114615: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18394;
 end   
18'd114616: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18394;
 end   
18'd114617: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18394;
 end   
18'd114618: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18394;
 end   
18'd114742: begin  
rid<=1;
end
18'd114743: begin  
end
18'd114744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd114745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd114746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd114747: begin  
rid<=0;
end
18'd114801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=69;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3584;
 end   
18'd114802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=47;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd114803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd114804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd114942: begin  
rid<=1;
end
18'd114943: begin  
end
18'd114944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd114945: begin  
rid<=0;
end
18'd115001: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=61;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5100;
 end   
18'd115002: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=20;
   mapp<=52;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5575;
 end   
18'd115003: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=80;
   mapp<=5;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=7202;
 end   
18'd115004: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=41;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=5285;
 end   
18'd115005: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=50;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=5258;
 end   
18'd115006: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=39;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=4486;
 end   
18'd115007: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=38;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=3843;
 end   
18'd115008: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=24;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=4187;
 end   
18'd115009: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=51;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd115010: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=5;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd115011: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd115012: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd115013: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5100;
 end   
18'd115142: begin  
rid<=1;
end
18'd115143: begin  
end
18'd115144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd115145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd115146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd115147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd115148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd115149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd115150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd115151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd115152: begin  
rid<=0;
end
18'd115201: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=4;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4446;
 end   
18'd115202: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=53;
   mapp<=82;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7895;
 end   
18'd115203: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=80;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=4480;
 end   
18'd115204: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=30;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=1682;
 end   
18'd115205: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=11;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=807;
 end   
18'd115206: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=6;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=4956;
 end   
18'd115207: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=58;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=8644;
 end   
18'd115208: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=87;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=6427;
 end   
18'd115209: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=51;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd115210: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd115211: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd115342: begin  
rid<=1;
end
18'd115343: begin  
end
18'd115344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd115345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd115346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd115347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd115348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd115349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd115350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd115351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd115352: begin  
rid<=0;
end
18'd115401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=96;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2770;
 end   
18'd115402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=14;
   mapp<=47;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4620;
 end   
18'd115403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd115404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd115405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd115542: begin  
rid<=1;
end
18'd115543: begin  
end
18'd115544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd115545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd115546: begin  
rid<=0;
end
18'd115601: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=10;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=60;
 end   
18'd115602: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=15;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=100;
 end   
18'd115603: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd115742: begin  
rid<=1;
end
18'd115743: begin  
end
18'd115744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd115745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd115746: begin  
rid<=0;
end
18'd115801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=13;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1887;
 end   
18'd115802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=23;
   mapp<=34;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4549;
 end   
18'd115803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=76;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8622;
 end   
18'd115804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=63;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=8003;
 end   
18'd115805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=77;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=7469;
 end   
18'd115806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=26;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=3008;
 end   
18'd115807: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=22;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=2168;
 end   
18'd115808: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=7;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd115809: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd115810: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd115942: begin  
rid<=1;
end
18'd115943: begin  
end
18'd115944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd115945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd115946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd115947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd115948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd115949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd115950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd115951: begin  
rid<=0;
end
18'd116001: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=25;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=675;
 end   
18'd116002: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10;
 end   
18'd116003: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=48;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1316;
 end   
18'd116004: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=75;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=2055;
 end   
18'd116005: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=30;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=850;
 end   
18'd116006: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd116142: begin  
rid<=1;
end
18'd116143: begin  
end
18'd116144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd116145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd116146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd116147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd116148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd116149: begin  
rid<=0;
end
18'd116201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=5;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1940;
 end   
18'd116202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=51;
   mapp<=16;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7778;
 end   
18'd116203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=7;
   mapp<=92;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1448;
 end   
18'd116204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=30;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=7282;
 end   
18'd116205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=3;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=5864;
 end   
18'd116206: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=47;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=10454;
 end   
18'd116207: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=52;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd116208: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=55;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd116209: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd116210: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd116211: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd116342: begin  
rid<=1;
end
18'd116343: begin  
end
18'd116344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd116345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd116346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd116347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd116348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd116349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd116350: begin  
rid<=0;
end
18'd116401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=99;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=36061;
 end   
18'd116402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=22;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd116403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=92;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd116404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=13;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd116405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=8;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd116406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=52;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd116407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=41;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd116408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=91;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd116409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=76;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd116410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=24;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd116411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=57;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd116412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd116413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=36061;
 end   
18'd116414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=36061;
 end   
18'd116415: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=36061;
 end   
18'd116416: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=36061;
 end   
18'd116417: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=36061;
 end   
18'd116418: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=36061;
 end   
18'd116419: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=36061;
 end   
18'd116420: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=36061;
 end   
18'd116421: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=36061;
 end   
18'd116422: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=36061;
 end   
18'd116542: begin  
rid<=1;
end
18'd116543: begin  
end
18'd116544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd116545: begin  
rid<=0;
end
18'd116601: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=9;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=20067;
 end   
18'd116602: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=50;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=21927;
 end   
18'd116603: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=54;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd116604: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=40;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd116605: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=97;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd116606: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=27;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd116607: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=79;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd116608: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=46;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd116609: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=39;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd116610: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=38;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd116611: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=81;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd116612: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd116613: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20067;
 end   
18'd116614: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20067;
 end   
18'd116615: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20067;
 end   
18'd116616: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20067;
 end   
18'd116617: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20067;
 end   
18'd116618: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20067;
 end   
18'd116619: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20067;
 end   
18'd116620: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20067;
 end   
18'd116621: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20067;
 end   
18'd116742: begin  
rid<=1;
end
18'd116743: begin  
end
18'd116744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd116745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd116746: begin  
rid<=0;
end
18'd116801: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=16;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14132;
 end   
18'd116802: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=94;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11326;
 end   
18'd116803: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=38;
   mapp<=93;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5510;
 end   
18'd116804: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=88;
   mapp<=13;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=10088;
 end   
18'd116805: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=6;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=10884;
 end   
18'd116806: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd116807: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd116808: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd116809: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd116810: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd116811: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd116812: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd116942: begin  
rid<=1;
end
18'd116943: begin  
end
18'd116944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd116945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd116946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd116947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd116948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd116949: begin  
rid<=0;
end
18'd117001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=56;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1896;
 end   
18'd117002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=9;
   mapp<=80;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5237;
 end   
18'd117003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=83;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=5262;
 end   
18'd117004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=66;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=4617;
 end   
18'd117005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd117006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd117007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd117142: begin  
rid<=1;
end
18'd117143: begin  
end
18'd117144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd117145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd117146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd117147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd117148: begin  
rid<=0;
end
18'd117201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=28;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13270;
 end   
18'd117202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=94;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=14140;
 end   
18'd117203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=32;
   mapp<=84;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=13050;
 end   
18'd117204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=66;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=14978;
 end   
18'd117205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=58;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=15024;
 end   
18'd117206: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=66;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=11021;
 end   
18'd117207: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=63;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd117208: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=13;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd117209: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd117210: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd117211: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd117342: begin  
rid<=1;
end
18'd117343: begin  
end
18'd117344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd117345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd117346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd117347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd117348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd117349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd117350: begin  
rid<=0;
end
18'd117401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=6;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=21584;
 end   
18'd117402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=46;
   mapp<=66;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=24290;
 end   
18'd117403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=74;
   mapp<=49;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=25645;
 end   
18'd117404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=8;
   mapp<=22;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=24579;
 end   
18'd117405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=46;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd117406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=70;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd117407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=20;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd117408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=66;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd117409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=69;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd117410: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=78;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd117411: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=27;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd117412: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd117413: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21584;
 end   
18'd117414: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21584;
 end   
18'd117415: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21584;
 end   
18'd117416: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21584;
 end   
18'd117417: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21584;
 end   
18'd117418: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21584;
 end   
18'd117419: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21584;
 end   
18'd117542: begin  
rid<=1;
end
18'd117543: begin  
end
18'd117544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd117545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd117546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd117547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd117548: begin  
rid<=0;
end
18'd117601: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=91;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=20162;
 end   
18'd117602: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=90;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=15400;
 end   
18'd117603: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=93;
   mapp<=78;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=10207;
 end   
18'd117604: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=44;
   mapp<=30;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=5458;
 end   
18'd117605: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=9;
   mapp<=21;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=5312;
 end   
18'd117606: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=7;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=6584;
 end   
18'd117607: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=40;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd117608: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd117609: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=22;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd117610: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=47;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd117611: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd117612: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd117613: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20162;
 end   
18'd117614: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20162;
 end   
18'd117615: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20162;
 end   
18'd117742: begin  
rid<=1;
end
18'd117743: begin  
end
18'd117744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd117745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd117746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd117747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd117748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd117749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd117750: begin  
rid<=0;
end
18'd117801: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=63;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10384;
 end   
18'd117802: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=79;
   mapp<=82;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10627;
 end   
18'd117803: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=69;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=7527;
 end   
18'd117804: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=40;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=2629;
 end   
18'd117805: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=1;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=4448;
 end   
18'd117806: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=55;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=3910;
 end   
18'd117807: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=5;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=2429;
 end   
18'd117808: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=26;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=8581;
 end   
18'd117809: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd117810: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd117811: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd117942: begin  
rid<=1;
end
18'd117943: begin  
end
18'd117944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd117945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd117946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd117947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd117948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd117949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd117950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd117951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd117952: begin  
rid<=0;
end
18'd118001: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=38;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10087;
 end   
18'd118002: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=17;
   mapp<=9;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2564;
 end   
18'd118003: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=95;
   mapp<=86;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5677;
 end   
18'd118004: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=9;
   mapp<=6;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=4737;
 end   
18'd118005: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=20;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=2479;
 end   
18'd118006: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=43;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=6325;
 end   
18'd118007: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=6;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=7544;
 end   
18'd118008: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd118009: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd118010: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd118011: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd118012: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd118013: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10087;
 end   
18'd118014: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10087;
 end   
18'd118142: begin  
rid<=1;
end
18'd118143: begin  
end
18'd118144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd118145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd118146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd118147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd118148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd118149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd118150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd118151: begin  
rid<=0;
end
18'd118201: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=62;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=21142;
 end   
18'd118202: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=97;
   mapp<=42;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=15038;
 end   
18'd118203: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=50;
   mapp<=52;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=15860;
 end   
18'd118204: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=89;
   mapp<=67;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=16944;
 end   
18'd118205: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=65;
   mapp<=40;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=14116;
 end   
18'd118206: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=5;
   mapp<=3;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=16814;
 end   
18'd118207: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd118208: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd118209: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd118210: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd118211: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd118212: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd118213: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21142;
 end   
18'd118214: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21142;
 end   
18'd118215: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21142;
 end   
18'd118216: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21142;
 end   
18'd118217: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21142;
 end   
18'd118342: begin  
rid<=1;
end
18'd118343: begin  
end
18'd118344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd118345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd118346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd118347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd118348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd118349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd118350: begin  
rid<=0;
end
18'd118401: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=60;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12829;
 end   
18'd118402: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=16;
   mapp<=3;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=12446;
 end   
18'd118403: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=81;
   mapp<=76;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=15237;
 end   
18'd118404: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=77;
   mapp<=65;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=15093;
 end   
18'd118405: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=75;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=12068;
 end   
18'd118406: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=46;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=5504;
 end   
18'd118407: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=81;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=11034;
 end   
18'd118408: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd118409: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd118410: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd118411: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd118412: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd118413: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12829;
 end   
18'd118414: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12829;
 end   
18'd118542: begin  
rid<=1;
end
18'd118543: begin  
end
18'd118544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd118545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd118546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd118547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd118548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd118549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd118550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd118551: begin  
rid<=0;
end
18'd118601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=2;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15495;
 end   
18'd118602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=35;
   mapp<=3;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11780;
 end   
18'd118603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=41;
   mapp<=44;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9745;
 end   
18'd118604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=86;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd118605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=93;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd118606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd118607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd118608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd118609: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd118610: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd118611: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd118612: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd118742: begin  
rid<=1;
end
18'd118743: begin  
end
18'd118744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd118745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd118746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd118747: begin  
rid<=0;
end
18'd118801: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=33;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11157;
 end   
18'd118802: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=11;
   mapp<=57;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13171;
 end   
18'd118803: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=76;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd118804: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=5;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd118805: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=65;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd118806: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=6;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd118807: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=98;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd118808: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=18;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd118809: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=19;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd118810: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd118811: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd118812: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd118813: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11157;
 end   
18'd118814: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11157;
 end   
18'd118815: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11157;
 end   
18'd118816: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11157;
 end   
18'd118817: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11157;
 end   
18'd118818: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11157;
 end   
18'd118819: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11157;
 end   
18'd118942: begin  
rid<=1;
end
18'd118943: begin  
end
18'd118944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd118945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd118946: begin  
rid<=0;
end
18'd119001: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=94;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=22273;
 end   
18'd119002: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=87;
   mapp<=50;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=20002;
 end   
18'd119003: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=65;
   mapp<=34;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=20211;
 end   
18'd119004: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=62;
   mapp<=95;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=24706;
 end   
18'd119005: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=39;
   mapp<=75;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=26458;
 end   
18'd119006: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=8;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd119007: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=60;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd119008: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=82;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd119009: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=86;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd119010: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=95;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd119011: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd119012: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd119013: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22273;
 end   
18'd119014: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22273;
 end   
18'd119015: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22273;
 end   
18'd119016: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22273;
 end   
18'd119142: begin  
rid<=1;
end
18'd119143: begin  
end
18'd119144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd119145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd119146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd119147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd119148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd119149: begin  
rid<=0;
end
18'd119201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=66;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10705;
 end   
18'd119202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=73;
   mapp<=59;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9162;
 end   
18'd119203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=50;
   mapp<=19;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=10273;
 end   
18'd119204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=60;
   mapp<=38;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=8920;
 end   
18'd119205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=41;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=8635;
 end   
18'd119206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=93;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=8144;
 end   
18'd119207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=48;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd119208: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=6;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd119209: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=18;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd119210: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd119211: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd119212: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd119213: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10705;
 end   
18'd119342: begin  
rid<=1;
end
18'd119343: begin  
end
18'd119344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd119345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd119346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd119347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd119348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd119349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd119350: begin  
rid<=0;
end
18'd119401: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=27;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3104;
 end   
18'd119402: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=71;
   mapp<=19;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4891;
 end   
18'd119403: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=14;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1728;
 end   
18'd119404: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=42;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd119405: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd119406: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd119542: begin  
rid<=1;
end
18'd119543: begin  
end
18'd119544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd119545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd119546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd119547: begin  
rid<=0;
end
18'd119601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=83;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5942;
 end   
18'd119602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=53;
   mapp<=61;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9334;
 end   
18'd119603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=5;
   mapp<=77;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8444;
 end   
18'd119604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=36;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=4373;
 end   
18'd119605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=25;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=2758;
 end   
18'd119606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd119607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd119608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd119609: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd119610: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd119742: begin  
rid<=1;
end
18'd119743: begin  
end
18'd119744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd119745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd119746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd119747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd119748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd119749: begin  
rid<=0;
end
18'd119801: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=44;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5065;
 end   
18'd119802: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=49;
   mapp<=45;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3313;
 end   
18'd119803: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=27;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=5128;
 end   
18'd119804: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=80;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=5069;
 end   
18'd119805: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=31;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=5324;
 end   
18'd119806: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=80;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=7637;
 end   
18'd119807: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=83;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=6015;
 end   
18'd119808: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=47;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=3265;
 end   
18'd119809: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=23;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=5061;
 end   
18'd119810: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=81;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[9]<=6741;
 end   
18'd119811: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd119812: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd119813: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5065;
 end   
18'd119942: begin  
rid<=1;
end
18'd119943: begin  
end
18'd119944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd119945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd119946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd119947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd119948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd119949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd119950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd119951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd119952: begin  
check<=expctdoutput[8]-outcheck;
end
18'd119953: begin  
check<=expctdoutput[9]-outcheck;
end
18'd119954: begin  
rid<=0;
end
18'd120001: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=27;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=22085;
 end   
18'd120002: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=25;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd120003: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=60;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd120004: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=69;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd120005: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=80;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd120006: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=23;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd120007: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd120008: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd120009: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd120010: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd120011: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd120012: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd120142: begin  
rid<=1;
end
18'd120143: begin  
end
18'd120144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd120145: begin  
rid<=0;
end
18'd120201: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=82;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5330;
 end   
18'd120202: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd120342: begin  
rid<=1;
end
18'd120343: begin  
end
18'd120344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd120345: begin  
rid<=0;
end
18'd120401: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=9;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=993;
 end   
18'd120402: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=30;
   mapp<=7;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3257;
 end   
18'd120403: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=91;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8014;
 end   
18'd120404: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=11;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=1295;
 end   
18'd120405: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=44;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=4176;
 end   
18'd120406: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=44;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=4403;
 end   
18'd120407: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=75;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=7208;
 end   
18'd120408: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=89;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=7848;
 end   
18'd120409: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=5;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd120410: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd120411: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd120542: begin  
rid<=1;
end
18'd120543: begin  
end
18'd120544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd120545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd120546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd120547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd120548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd120549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd120550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd120551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd120552: begin  
rid<=0;
end
18'd120601: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=50;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=19206;
 end   
18'd120602: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=88;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=18938;
 end   
18'd120603: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=66;
   mapp<=48;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=16458;
 end   
18'd120604: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=67;
   mapp<=60;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=15461;
 end   
18'd120605: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=78;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd120606: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=73;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd120607: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=43;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd120608: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=48;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd120609: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd120610: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd120611: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd120612: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd120613: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19206;
 end   
18'd120742: begin  
rid<=1;
end
18'd120743: begin  
end
18'd120744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd120745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd120746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd120747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd120748: begin  
rid<=0;
end
18'd120801: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=57;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14717;
 end   
18'd120802: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=80;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd120803: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=66;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd120804: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=61;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd120805: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd120806: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd120807: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd120808: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd120942: begin  
rid<=1;
end
18'd120943: begin  
end
18'd120944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd120945: begin  
rid<=0;
end
18'd121001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=88;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=25006;
 end   
18'd121002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=88;
   mapp<=85;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=20602;
 end   
18'd121003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=86;
   mapp<=50;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=13696;
 end   
18'd121004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=57;
   mapp<=91;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=11376;
 end   
18'd121005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=59;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd121006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=27;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd121007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=10;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd121008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=26;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd121009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd121010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd121011: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd121012: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd121013: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25006;
 end   
18'd121142: begin  
rid<=1;
end
18'd121143: begin  
end
18'd121144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd121145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd121146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd121147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd121148: begin  
rid<=0;
end
18'd121201: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=92;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5888;
 end   
18'd121202: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=66;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=6082;
 end   
18'd121203: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=74;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=6828;
 end   
18'd121204: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=92;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=8494;
 end   
18'd121205: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=48;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=4456;
 end   
18'd121206: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=12;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=1154;
 end   
18'd121207: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd121342: begin  
rid<=1;
end
18'd121343: begin  
end
18'd121344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd121345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd121346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd121347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd121348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd121349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd121350: begin  
rid<=0;
end
18'd121401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=96;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=19326;
 end   
18'd121402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=96;
   mapp<=59;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=21082;
 end   
18'd121403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=78;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd121404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=8;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd121405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=86;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd121406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=37;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd121407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=3;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd121408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd121409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd121410: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd121411: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd121412: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd121413: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19326;
 end   
18'd121414: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19326;
 end   
18'd121415: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19326;
 end   
18'd121542: begin  
rid<=1;
end
18'd121543: begin  
end
18'd121544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd121545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd121546: begin  
rid<=0;
end
18'd121601: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=4;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13259;
 end   
18'd121602: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=42;
   mapp<=45;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13561;
 end   
18'd121603: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=24;
   mapp<=30;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=18921;
 end   
18'd121604: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=69;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd121605: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=81;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd121606: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=43;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd121607: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd121608: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd121609: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd121610: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd121611: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd121612: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd121613: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13259;
 end   
18'd121614: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13259;
 end   
18'd121742: begin  
rid<=1;
end
18'd121743: begin  
end
18'd121744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd121745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd121746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd121747: begin  
rid<=0;
end
18'd121801: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=34;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=281;
 end   
18'd121802: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=1;
   mapp<=23;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2079;
 end   
18'd121803: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=5;
   mapp<=38;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=4662;
 end   
18'd121804: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=61;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=5090;
 end   
18'd121805: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=32;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=3370;
 end   
18'd121806: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=56;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd121807: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=36;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd121808: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=10;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd121809: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd121810: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd121811: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd121812: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd121942: begin  
rid<=1;
end
18'd121943: begin  
end
18'd121944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd121945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd121946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd121947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd121948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd121949: begin  
rid<=0;
end
18'd122001: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=90;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8416;
 end   
18'd122002: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=8;
   mapp<=92;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8416;
 end   
18'd122003: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=75;
   mapp<=10;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=14673;
 end   
18'd122004: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=89;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=14141;
 end   
18'd122005: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=69;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=14115;
 end   
18'd122006: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=91;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=10995;
 end   
18'd122007: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=39;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=6343;
 end   
18'd122008: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=35;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=3707;
 end   
18'd122009: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=6;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd122010: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=39;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd122011: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd122012: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd122013: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8416;
 end   
18'd122142: begin  
rid<=1;
end
18'd122143: begin  
end
18'd122144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd122145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd122146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd122147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd122148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd122149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd122150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd122151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd122152: begin  
rid<=0;
end
18'd122201: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=64;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14128;
 end   
18'd122202: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=48;
   mapp<=44;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8234;
 end   
18'd122203: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=8;
   mapp<=27;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=13452;
 end   
18'd122204: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=72;
   mapp<=95;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=8870;
 end   
18'd122205: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=8;
   mapp<=36;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=8128;
 end   
18'd122206: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=95;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=7034;
 end   
18'd122207: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd122208: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd122209: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd122210: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd122211: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd122212: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd122213: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14128;
 end   
18'd122214: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14128;
 end   
18'd122215: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14128;
 end   
18'd122342: begin  
rid<=1;
end
18'd122343: begin  
end
18'd122344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd122345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd122346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd122347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd122348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd122349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd122350: begin  
rid<=0;
end
18'd122401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=67;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=19293;
 end   
18'd122402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=5;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd122403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=11;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd122404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=83;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd122405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=53;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd122406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=39;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd122407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=26;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd122408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=42;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd122409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd122410: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd122411: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd122412: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd122413: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19293;
 end   
18'd122414: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19293;
 end   
18'd122415: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19293;
 end   
18'd122416: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19293;
 end   
18'd122542: begin  
rid<=1;
end
18'd122543: begin  
end
18'd122544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd122545: begin  
rid<=0;
end
18'd122601: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=70;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6444;
 end   
18'd122602: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=10;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8071;
 end   
18'd122603: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=5;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd122604: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=9;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd122605: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=71;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd122606: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd122607: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd122608: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd122609: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd122610: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd122611: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd122742: begin  
rid<=1;
end
18'd122743: begin  
end
18'd122744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd122745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd122746: begin  
rid<=0;
end
18'd122801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=88;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12688;
 end   
18'd122802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=51;
   mapp<=42;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11813;
 end   
18'd122803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=52;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd122804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=57;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd122805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=65;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd122806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd122807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd122808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd122809: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd122810: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd122811: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd122942: begin  
rid<=1;
end
18'd122943: begin  
end
18'd122944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd122945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd122946: begin  
rid<=0;
end
18'd123001: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=60;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=28710;
 end   
18'd123002: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=56;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=27577;
 end   
18'd123003: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=92;
   mapp<=50;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=36108;
 end   
18'd123004: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=93;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd123005: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=99;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd123006: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=32;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd123007: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=49;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd123008: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=73;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd123009: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd123010: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd123011: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd123012: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd123013: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28710;
 end   
18'd123014: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28710;
 end   
18'd123015: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28710;
 end   
18'd123016: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28710;
 end   
18'd123017: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28710;
 end   
18'd123018: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=28710;
 end   
18'd123142: begin  
rid<=1;
end
18'd123143: begin  
end
18'd123144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd123145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd123146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd123147: begin  
rid<=0;
end
18'd123201: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=9;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9758;
 end   
18'd123202: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=95;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9859;
 end   
18'd123203: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=47;
   mapp<=86;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6177;
 end   
18'd123204: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=25;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=6335;
 end   
18'd123205: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=64;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=2120;
 end   
18'd123206: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=4124;
 end   
18'd123207: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=32;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=4553;
 end   
18'd123208: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=22;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=7034;
 end   
18'd123209: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd123210: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd123211: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd123212: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd123213: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9758;
 end   
18'd123342: begin  
rid<=1;
end
18'd123343: begin  
end
18'd123344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd123345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd123346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd123347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd123348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd123349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd123350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd123351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd123352: begin  
rid<=0;
end
18'd123401: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=65;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6006;
 end   
18'd123402: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=62;
   mapp<=36;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6768;
 end   
18'd123403: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=68;
   mapp<=23;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9819;
 end   
18'd123404: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=44;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=14094;
 end   
18'd123405: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=82;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=16050;
 end   
18'd123406: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=90;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=13678;
 end   
18'd123407: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=75;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=10439;
 end   
18'd123408: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=46;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=8742;
 end   
18'd123409: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd123410: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd123411: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd123412: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd123413: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6006;
 end   
18'd123542: begin  
rid<=1;
end
18'd123543: begin  
end
18'd123544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd123545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd123546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd123547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd123548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd123549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd123550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd123551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd123552: begin  
rid<=0;
end
18'd123601: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=87;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7654;
 end   
18'd123602: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=40;
   mapp<=13;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4148;
 end   
18'd123603: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=66;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5861;
 end   
18'd123604: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=33;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd123605: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd123606: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd123742: begin  
rid<=1;
end
18'd123743: begin  
end
18'd123744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd123745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd123746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd123747: begin  
rid<=0;
end
18'd123801: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=33;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16169;
 end   
18'd123802: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=66;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=15047;
 end   
18'd123803: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=55;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd123804: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=57;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd123805: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=21;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd123806: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=61;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd123807: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=1;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd123808: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd123809: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd123810: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd123811: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd123812: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd123813: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16169;
 end   
18'd123814: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16169;
 end   
18'd123815: begin  
  clrr<=0;
  maplen<=8;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16169;
 end   
18'd123942: begin  
rid<=1;
end
18'd123943: begin  
end
18'd123944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd123945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd123946: begin  
rid<=0;
end
18'd124001: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=99;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=36172;
 end   
18'd124002: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=15;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd124003: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=66;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd124004: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=65;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd124005: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=32;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd124006: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=74;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd124007: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=78;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd124008: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=37;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd124009: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd124010: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd124011: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd124012: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd124013: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=36172;
 end   
18'd124014: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=36172;
 end   
18'd124015: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=36172;
 end   
18'd124016: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=36172;
 end   
18'd124142: begin  
rid<=1;
end
18'd124143: begin  
end
18'd124144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd124145: begin  
rid<=0;
end
18'd124201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=58;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5394;
 end   
18'd124202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=58;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=3374;
 end   
18'd124203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=57;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=3326;
 end   
18'd124204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=71;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=4148;
 end   
18'd124205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd124342: begin  
rid<=1;
end
18'd124343: begin  
end
18'd124344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd124345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd124346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd124347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd124348: begin  
rid<=0;
end
18'd124401: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=78;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15857;
 end   
18'd124402: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=6;
   mapp<=6;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11572;
 end   
18'd124403: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=24;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd124404: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=15;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd124405: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=73;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd124406: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=60;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd124407: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=78;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd124408: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=36;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd124409: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=19;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd124410: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd124411: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd124412: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd124413: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15857;
 end   
18'd124414: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15857;
 end   
18'd124415: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15857;
 end   
18'd124416: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15857;
 end   
18'd124417: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15857;
 end   
18'd124418: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15857;
 end   
18'd124419: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15857;
 end   
18'd124542: begin  
rid<=1;
end
18'd124543: begin  
end
18'd124544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd124545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd124546: begin  
rid<=0;
end
18'd124601: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=16;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1795;
 end   
18'd124602: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=23;
   mapp<=21;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2148;
 end   
18'd124603: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=12;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=2810;
 end   
18'd124604: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=86;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=8552;
 end   
18'd124605: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=70;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=7166;
 end   
18'd124606: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=66;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=6344;
 end   
18'd124607: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=42;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=4932;
 end   
18'd124608: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=68;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=6864;
 end   
18'd124609: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=58;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=6432;
 end   
18'd124610: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=76;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd124611: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd124612: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd124742: begin  
rid<=1;
end
18'd124743: begin  
end
18'd124744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd124745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd124746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd124747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd124748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd124749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd124750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd124751: begin  
check<=expctdoutput[7]-outcheck;
end
18'd124752: begin  
check<=expctdoutput[8]-outcheck;
end
18'd124753: begin  
rid<=0;
end
18'd124801: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=21;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6642;
 end   
18'd124802: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=37;
   mapp<=53;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8989;
 end   
18'd124803: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=4;
   mapp<=4;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=3614;
 end   
18'd124804: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=78;
   mapp<=38;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=11915;
 end   
18'd124805: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=97;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=4129;
 end   
18'd124806: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=22;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=5241;
 end   
18'd124807: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=95;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=9308;
 end   
18'd124808: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd124809: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd124810: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd124811: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd124812: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd124813: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6642;
 end   
18'd124814: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6642;
 end   
18'd124942: begin  
rid<=1;
end
18'd124943: begin  
end
18'd124944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd124945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd124946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd124947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd124948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd124949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd124950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd124951: begin  
rid<=0;
end
18'd125001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=89;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11088;
 end   
18'd125002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=2;
   mapp<=94;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13388;
 end   
18'd125003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=11;
   mapp<=31;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8810;
 end   
18'd125004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=57;
   mapp<=65;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=11053;
 end   
18'd125005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=7;
   mapp<=56;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=6704;
 end   
18'd125006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=7;
   mapp<=84;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=12015;
 end   
18'd125007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd125008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd125009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd125010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd125011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd125012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd125013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11088;
 end   
18'd125014: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11088;
 end   
18'd125015: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11088;
 end   
18'd125016: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11088;
 end   
18'd125017: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11088;
 end   
18'd125142: begin  
rid<=1;
end
18'd125143: begin  
end
18'd125144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd125145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd125146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd125147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd125148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd125149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd125150: begin  
rid<=0;
end
18'd125201: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=35;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3823;
 end   
18'd125202: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=46;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3616;
 end   
18'd125203: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=59;
   mapp<=12;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6409;
 end   
18'd125204: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=31;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=7548;
 end   
18'd125205: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=77;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=5343;
 end   
18'd125206: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=49;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=2100;
 end   
18'd125207: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd125208: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd125209: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd125210: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd125211: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd125342: begin  
rid<=1;
end
18'd125343: begin  
end
18'd125344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd125345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd125346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd125347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd125348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd125349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd125350: begin  
rid<=0;
end
18'd125401: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=80;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13240;
 end   
18'd125402: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=55;
   mapp<=90;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=18176;
 end   
18'd125403: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=68;
   mapp<=64;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12413;
 end   
18'd125404: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=34;
   mapp<=97;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=12463;
 end   
18'd125405: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=25;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=8579;
 end   
18'd125406: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=7;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=8813;
 end   
18'd125407: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=83;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=15957;
 end   
18'd125408: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd125409: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd125410: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd125411: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd125412: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd125413: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13240;
 end   
18'd125414: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13240;
 end   
18'd125542: begin  
rid<=1;
end
18'd125543: begin  
end
18'd125544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd125545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd125546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd125547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd125548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd125549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd125550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd125551: begin  
rid<=0;
end
18'd125601: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=23;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=21620;
 end   
18'd125602: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=87;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd125603: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=78;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd125604: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=39;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd125605: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=3;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd125606: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=37;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd125607: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=90;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd125608: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=63;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd125609: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=77;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd125610: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=1;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd125611: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd125612: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd125613: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21620;
 end   
18'd125614: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21620;
 end   
18'd125615: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21620;
 end   
18'd125616: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21620;
 end   
18'd125617: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21620;
 end   
18'd125618: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21620;
 end   
18'd125619: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21620;
 end   
18'd125620: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21620;
 end   
18'd125742: begin  
rid<=1;
end
18'd125743: begin  
end
18'd125744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd125745: begin  
rid<=0;
end
18'd125801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=90;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3652;
 end   
18'd125802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=68;
   mapp<=14;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8002;
 end   
18'd125803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=99;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=15594;
 end   
18'd125804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=98;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=9054;
 end   
18'd125805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=3;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=6974;
 end   
18'd125806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=98;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=10026;
 end   
18'd125807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd125808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd125809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd125942: begin  
rid<=1;
end
18'd125943: begin  
end
18'd125944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd125945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd125946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd125947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd125948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd125949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd125950: begin  
rid<=0;
end
18'd126001: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=35;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13738;
 end   
18'd126002: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=7;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd126003: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=77;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd126004: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=71;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd126005: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=5;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd126006: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=30;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd126007: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd126008: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd126009: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd126010: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd126011: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd126012: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd126142: begin  
rid<=1;
end
18'd126143: begin  
end
18'd126144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd126145: begin  
rid<=0;
end
18'd126201: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=59;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3422;
 end   
18'd126202: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=98;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5694;
 end   
18'd126203: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=42;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=2456;
 end   
18'd126204: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=8;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=494;
 end   
18'd126205: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=77;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=4506;
 end   
18'd126206: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd126342: begin  
rid<=1;
end
18'd126343: begin  
end
18'd126344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd126345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd126346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd126347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd126348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd126349: begin  
rid<=0;
end
18'd126401: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=26;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4810;
 end   
18'd126402: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=60;
   mapp<=78;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7438;
 end   
18'd126403: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=90;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=3020;
 end   
18'd126404: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=11;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=2716;
 end   
18'd126405: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=40;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=2100;
 end   
18'd126406: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=17;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=612;
 end   
18'd126407: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=2;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=4252;
 end   
18'd126408: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=69;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=4444;
 end   
18'd126409: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=43;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=4078;
 end   
18'd126410: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd126411: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd126412: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd126542: begin  
rid<=1;
end
18'd126543: begin  
end
18'd126544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd126545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd126546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd126547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd126548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd126549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd126550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd126551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd126552: begin  
check<=expctdoutput[8]-outcheck;
end
18'd126553: begin  
rid<=0;
end
18'd126601: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=10;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13192;
 end   
18'd126602: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=49;
   mapp<=90;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13258;
 end   
18'd126603: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=39;
   mapp<=68;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=10428;
 end   
18'd126604: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=13;
   mapp<=26;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=13854;
 end   
18'd126605: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=62;
   mapp<=86;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=11724;
 end   
18'd126606: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=58;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=13874;
 end   
18'd126607: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=20;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd126608: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd126609: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=15;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd126610: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=75;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd126611: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd126612: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd126613: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13192;
 end   
18'd126614: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13192;
 end   
18'd126615: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13192;
 end   
18'd126742: begin  
rid<=1;
end
18'd126743: begin  
end
18'd126744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd126745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd126746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd126747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd126748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd126749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd126750: begin  
rid<=0;
end
18'd126801: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=77;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13841;
 end   
18'd126802: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=84;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd126803: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=75;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd126804: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=35;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd126805: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd126806: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd126807: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd126808: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd126942: begin  
rid<=1;
end
18'd126943: begin  
end
18'd126944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd126945: begin  
rid<=0;
end
18'd127001: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=23;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2409;
 end   
18'd127002: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=45;
   mapp<=29;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4727;
 end   
18'd127003: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=90;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=3575;
 end   
18'd127004: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=33;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=3804;
 end   
18'd127005: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=67;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=3246;
 end   
18'd127006: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd127007: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd127008: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd127142: begin  
rid<=1;
end
18'd127143: begin  
end
18'd127144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd127145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd127146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd127147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd127148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd127149: begin  
rid<=0;
end
18'd127201: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=4;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14689;
 end   
18'd127202: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=78;
   mapp<=34;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=22678;
 end   
18'd127203: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=91;
   mapp<=52;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=20639;
 end   
18'd127204: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=33;
   mapp<=75;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=11907;
 end   
18'd127205: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=60;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd127206: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=25;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd127207: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=26;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd127208: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=25;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd127209: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=90;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd127210: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd127211: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=7;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd127212: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd127213: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14689;
 end   
18'd127214: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14689;
 end   
18'd127215: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14689;
 end   
18'd127216: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14689;
 end   
18'd127217: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14689;
 end   
18'd127218: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14689;
 end   
18'd127219: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14689;
 end   
18'd127342: begin  
rid<=1;
end
18'd127343: begin  
end
18'd127344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd127345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd127346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd127347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd127348: begin  
rid<=0;
end
18'd127401: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=9;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=18421;
 end   
18'd127402: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=66;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd127403: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=65;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd127404: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=65;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd127405: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=87;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd127406: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=73;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd127407: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=76;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd127408: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=50;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd127409: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=53;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd127410: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd127411: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd127412: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd127413: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18421;
 end   
18'd127414: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18421;
 end   
18'd127415: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18421;
 end   
18'd127416: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18421;
 end   
18'd127417: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18421;
 end   
18'd127418: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18421;
 end   
18'd127542: begin  
rid<=1;
end
18'd127543: begin  
end
18'd127544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd127545: begin  
rid<=0;
end
18'd127601: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=68;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11477;
 end   
18'd127602: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=2;
   mapp<=43;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=17794;
 end   
18'd127603: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=60;
   mapp<=0;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=16533;
 end   
18'd127604: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=68;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd127605: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=73;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd127606: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=66;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd127607: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd127608: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd127609: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd127610: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd127611: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd127612: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd127613: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11477;
 end   
18'd127614: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11477;
 end   
18'd127742: begin  
rid<=1;
end
18'd127743: begin  
end
18'd127744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd127745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd127746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd127747: begin  
rid<=0;
end
18'd127801: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=94;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7990;
 end   
18'd127802: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=1;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=104;
 end   
18'd127803: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=85;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=8010;
 end   
18'd127804: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=19;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=1816;
 end   
18'd127805: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=46;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=4364;
 end   
18'd127806: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=13;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=1272;
 end   
18'd127807: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=96;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=9084;
 end   
18'd127808: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=89;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=8436;
 end   
18'd127809: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd127942: begin  
rid<=1;
end
18'd127943: begin  
end
18'd127944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd127945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd127946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd127947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd127948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd127949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd127950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd127951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd127952: begin  
rid<=0;
end
18'd128001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=52;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=988;
 end   
18'd128002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=27;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=1414;
 end   
18'd128003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=88;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=4596;
 end   
18'd128004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=61;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=3202;
 end   
18'd128005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=95;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=4980;
 end   
18'd128006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd128142: begin  
rid<=1;
end
18'd128143: begin  
end
18'd128144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd128145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd128146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd128147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd128148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd128149: begin  
rid<=0;
end
18'd128201: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=53;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8711;
 end   
18'd128202: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=92;
   mapp<=65;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6503;
 end   
18'd128203: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=10;
   mapp<=24;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9270;
 end   
18'd128204: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd128205: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd128206: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd128207: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd128208: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd128342: begin  
rid<=1;
end
18'd128343: begin  
end
18'd128344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd128345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd128346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd128347: begin  
rid<=0;
end
18'd128401: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=56;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3076;
 end   
18'd128402: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=65;
   mapp<=12;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6338;
 end   
18'd128403: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=36;
   mapp<=56;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=7876;
 end   
18'd128404: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=56;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=6232;
 end   
18'd128405: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=30;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=4959;
 end   
18'd128406: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=31;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=4032;
 end   
18'd128407: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=34;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=4585;
 end   
18'd128408: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=1;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=6109;
 end   
18'd128409: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd128410: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd128411: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd128412: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd128413: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=3076;
 end   
18'd128542: begin  
rid<=1;
end
18'd128543: begin  
end
18'd128544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd128545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd128546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd128547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd128548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd128549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd128550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd128551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd128552: begin  
rid<=0;
end
18'd128601: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=2;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3916;
 end   
18'd128602: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=52;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9594;
 end   
18'd128603: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=71;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=11886;
 end   
18'd128604: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=80;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd128605: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd128606: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd128742: begin  
rid<=1;
end
18'd128743: begin  
end
18'd128744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd128745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd128746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd128747: begin  
rid<=0;
end
18'd128801: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=67;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3752;
 end   
18'd128802: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=28;
   mapp<=99;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2569;
 end   
18'd128803: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=12;
   mapp<=37;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6293;
 end   
18'd128804: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=31;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=12035;
 end   
18'd128805: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=84;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=12065;
 end   
18'd128806: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=93;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=8016;
 end   
18'd128807: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=58;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=7703;
 end   
18'd128808: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=40;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd128809: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=87;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd128810: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd128811: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd128812: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd128942: begin  
rid<=1;
end
18'd128943: begin  
end
18'd128944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd128945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd128946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd128947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd128948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd128949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd128950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd128951: begin  
rid<=0;
end
18'd129001: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=60;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3540;
 end   
18'd129002: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=59;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=3550;
 end   
18'd129003: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=30;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=1820;
 end   
18'd129004: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=30;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=1830;
 end   
18'd129005: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=76;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=4600;
 end   
18'd129006: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=40;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=2450;
 end   
18'd129007: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=38;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=2340;
 end   
18'd129008: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=91;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=5530;
 end   
18'd129009: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=60;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=3680;
 end   
18'd129010: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=76;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[9]<=4650;
 end   
18'd129011: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd129142: begin  
rid<=1;
end
18'd129143: begin  
end
18'd129144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd129145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd129146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd129147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd129148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd129149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd129150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd129151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd129152: begin  
check<=expctdoutput[8]-outcheck;
end
18'd129153: begin  
check<=expctdoutput[9]-outcheck;
end
18'd129154: begin  
rid<=0;
end
18'd129201: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=28;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11708;
 end   
18'd129202: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=96;
   mapp<=53;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=15323;
 end   
18'd129203: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=4;
   mapp<=85;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=15208;
 end   
18'd129204: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=68;
   mapp<=39;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=16757;
 end   
18'd129205: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=96;
   mapp<=27;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=14366;
 end   
18'd129206: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=75;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd129207: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=13;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd129208: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=83;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd129209: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=91;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd129210: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd129211: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd129212: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd129213: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11708;
 end   
18'd129214: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11708;
 end   
18'd129342: begin  
rid<=1;
end
18'd129343: begin  
end
18'd129344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd129345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd129346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd129347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd129348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd129349: begin  
rid<=0;
end
18'd129401: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=95;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12077;
 end   
18'd129402: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=52;
   mapp<=59;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9943;
 end   
18'd129403: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=35;
   mapp<=27;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=11537;
 end   
18'd129404: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=60;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd129405: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=52;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd129406: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=71;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd129407: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=95;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd129408: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=20;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd129409: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd129410: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd129411: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd129412: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd129413: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12077;
 end   
18'd129414: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12077;
 end   
18'd129542: begin  
rid<=1;
end
18'd129543: begin  
end
18'd129544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd129545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd129546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd129547: begin  
rid<=0;
end
18'd129601: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=12;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9441;
 end   
18'd129602: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=74;
   mapp<=75;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10533;
 end   
18'd129603: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=49;
   mapp<=63;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=7317;
 end   
18'd129604: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=30;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=10125;
 end   
18'd129605: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=28;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=14270;
 end   
18'd129606: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=95;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd129607: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=83;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd129608: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd129609: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd129610: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd129742: begin  
rid<=1;
end
18'd129743: begin  
end
18'd129744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd129745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd129746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd129747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd129748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd129749: begin  
rid<=0;
end
18'd129801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=93;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15880;
 end   
18'd129802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=96;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=19132;
 end   
18'd129803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=73;
   mapp<=85;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=24139;
 end   
18'd129804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=61;
   mapp<=90;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=22417;
 end   
18'd129805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd129806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd129807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd129808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd129809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd129810: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd129811: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd129942: begin  
rid<=1;
end
18'd129943: begin  
end
18'd129944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd129945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd129946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd129947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd129948: begin  
rid<=0;
end
18'd130001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=78;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=18612;
 end   
18'd130002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=89;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd130003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=72;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd130004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=93;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd130005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=58;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd130006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd130007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd130008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd130009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd130010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd130142: begin  
rid<=1;
end
18'd130143: begin  
end
18'd130144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd130145: begin  
rid<=0;
end
18'd130201: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=2;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=31579;
 end   
18'd130202: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=26;
   mapp<=10;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=34843;
 end   
18'd130203: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=94;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd130204: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=45;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd130205: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=74;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd130206: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=48;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd130207: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=83;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd130208: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=44;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd130209: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=81;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd130210: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=75;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd130211: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd130212: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd130213: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=31579;
 end   
18'd130214: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=31579;
 end   
18'd130215: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=31579;
 end   
18'd130216: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=31579;
 end   
18'd130217: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=31579;
 end   
18'd130218: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=31579;
 end   
18'd130219: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=31579;
 end   
18'd130342: begin  
rid<=1;
end
18'd130343: begin  
end
18'd130344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd130345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd130346: begin  
rid<=0;
end
18'd130401: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=91;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=21420;
 end   
18'd130402: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=89;
   mapp<=98;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=26407;
 end   
18'd130403: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=68;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd130404: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=60;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd130405: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=12;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd130406: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd130407: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd130408: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd130409: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd130410: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd130411: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd130412: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd130413: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21420;
 end   
18'd130542: begin  
rid<=1;
end
18'd130543: begin  
end
18'd130544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd130545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd130546: begin  
rid<=0;
end
18'd130601: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=90;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=19596;
 end   
18'd130602: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=40;
   mapp<=75;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9421;
 end   
18'd130603: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=5;
   mapp<=17;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=11704;
 end   
18'd130604: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=84;
   mapp<=90;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=15721;
 end   
18'd130605: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=43;
   mapp<=47;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=10095;
 end   
18'd130606: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=14;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd130607: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=64;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd130608: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd130609: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=98;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd130610: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd130611: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd130612: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd130613: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19596;
 end   
18'd130614: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19596;
 end   
18'd130742: begin  
rid<=1;
end
18'd130743: begin  
end
18'd130744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd130745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd130746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd130747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd130748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd130749: begin  
rid<=0;
end
18'd130801: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=77;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16151;
 end   
18'd130802: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=23;
   mapp<=23;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=14427;
 end   
18'd130803: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=60;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd130804: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=64;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd130805: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=17;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd130806: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=67;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd130807: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd130808: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd130809: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd130810: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd130811: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd130942: begin  
rid<=1;
end
18'd130943: begin  
end
18'd130944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd130945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd130946: begin  
rid<=0;
end
18'd131001: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=65;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5951;
 end   
18'd131002: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10409;
 end   
18'd131003: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=88;
   mapp<=27;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=11904;
 end   
18'd131004: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=69;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=7732;
 end   
18'd131005: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=13;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd131006: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=98;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd131007: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd131008: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd131009: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd131142: begin  
rid<=1;
end
18'd131143: begin  
end
18'd131144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd131145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd131146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd131147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd131148: begin  
rid<=0;
end
18'd131201: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=5;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=810;
 end   
18'd131202: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=10;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2078;
 end   
18'd131203: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=28;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=2148;
 end   
18'd131204: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=13;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=1800;
 end   
18'd131205: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=20;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=5632;
 end   
18'd131206: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=82;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=5942;
 end   
18'd131207: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=32;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=5356;
 end   
18'd131208: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=66;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=8242;
 end   
18'd131209: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=87;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=6166;
 end   
18'd131210: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=31;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd131211: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd131212: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd131342: begin  
rid<=1;
end
18'd131343: begin  
end
18'd131344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd131345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd131346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd131347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd131348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd131349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd131350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd131351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd131352: begin  
check<=expctdoutput[8]-outcheck;
end
18'd131353: begin  
rid<=0;
end
18'd131401: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=94;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14039;
 end   
18'd131402: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=27;
   mapp<=85;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13402;
 end   
18'd131403: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=88;
   mapp<=2;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=20076;
 end   
18'd131404: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=54;
   mapp<=73;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=12107;
 end   
18'd131405: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=2;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd131406: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=66;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd131407: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=68;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd131408: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=47;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd131409: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd131410: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd131411: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd131412: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd131413: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14039;
 end   
18'd131542: begin  
rid<=1;
end
18'd131543: begin  
end
18'd131544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd131545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd131546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd131547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd131548: begin  
rid<=0;
end
18'd131601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=41;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5792;
 end   
18'd131602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=63;
   mapp<=12;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9085;
 end   
18'd131603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=48;
   mapp<=62;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=11325;
 end   
18'd131604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=32;
   mapp<=20;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=12035;
 end   
18'd131605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=67;
   mapp<=1;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=11517;
 end   
18'd131606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd131607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd131608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd131609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd131610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd131611: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd131612: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd131613: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5792;
 end   
18'd131614: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5792;
 end   
18'd131742: begin  
rid<=1;
end
18'd131743: begin  
end
18'd131744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd131745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd131746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd131747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd131748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd131749: begin  
rid<=0;
end
18'd131801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=7;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7141;
 end   
18'd131802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=75;
   mapp<=94;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7189;
 end   
18'd131803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=66;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=3604;
 end   
18'd131804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=29;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=8115;
 end   
18'd131805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=82;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=1858;
 end   
18'd131806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=8;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd131807: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd131808: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd131942: begin  
rid<=1;
end
18'd131943: begin  
end
18'd131944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd131945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd131946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd131947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd131948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd131949: begin  
rid<=0;
end
18'd132001: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=40;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=21602;
 end   
18'd132002: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=3;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd132003: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=25;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd132004: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=28;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd132005: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=59;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd132006: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=89;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd132007: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=70;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd132008: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=49;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd132009: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=12;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd132010: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=88;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd132011: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd132012: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd132013: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21602;
 end   
18'd132014: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21602;
 end   
18'd132015: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21602;
 end   
18'd132016: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21602;
 end   
18'd132017: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21602;
 end   
18'd132018: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21602;
 end   
18'd132019: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21602;
 end   
18'd132020: begin  
  clrr<=0;
  maplen<=10;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21602;
 end   
18'd132142: begin  
rid<=1;
end
18'd132143: begin  
end
18'd132144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd132145: begin  
rid<=0;
end
18'd132201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=11;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2185;
 end   
18'd132202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=75;
   mapp<=14;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6843;
 end   
18'd132203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=84;
   mapp<=5;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8106;
 end   
18'd132204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=6;
   mapp<=44;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=5709;
 end   
18'd132205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=58;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=6842;
 end   
18'd132206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=97;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd132207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=94;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd132208: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=59;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd132209: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd132210: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd132211: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd132212: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd132342: begin  
rid<=1;
end
18'd132343: begin  
end
18'd132344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd132345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd132346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd132347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd132348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd132349: begin  
rid<=0;
end
18'd132401: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=87;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=25777;
 end   
18'd132402: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=43;
   mapp<=22;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=26282;
 end   
18'd132403: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=41;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd132404: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=39;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd132405: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=88;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd132406: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=39;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd132407: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=77;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd132408: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=72;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd132409: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd132410: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd132411: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd132412: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd132413: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25777;
 end   
18'd132414: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25777;
 end   
18'd132415: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25777;
 end   
18'd132416: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25777;
 end   
18'd132417: begin  
  clrr<=0;
  maplen<=9;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25777;
 end   
18'd132542: begin  
rid<=1;
end
18'd132543: begin  
end
18'd132544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd132545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd132546: begin  
rid<=0;
end
18'd132601: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=99;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=17588;
 end   
18'd132602: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=15;
   mapp<=71;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=14135;
 end   
18'd132603: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=22;
   mapp<=85;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=17330;
 end   
18'd132604: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=42;
   mapp<=29;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=20728;
 end   
18'd132605: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=12;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd132606: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=7;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd132607: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=31;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd132608: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=48;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd132609: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=54;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd132610: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=71;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd132611: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=90;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd132612: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd132613: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17588;
 end   
18'd132614: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17588;
 end   
18'd132615: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17588;
 end   
18'd132616: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17588;
 end   
18'd132617: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17588;
 end   
18'd132618: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17588;
 end   
18'd132619: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17588;
 end   
18'd132742: begin  
rid<=1;
end
18'd132743: begin  
end
18'd132744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd132745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd132746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd132747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd132748: begin  
rid<=0;
end
18'd132801: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=23;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11810;
 end   
18'd132802: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=41;
   mapp<=27;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8845;
 end   
18'd132803: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=49;
   mapp<=68;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=14549;
 end   
18'd132804: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=34;
   mapp<=64;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=7616;
 end   
18'd132805: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=84;
   mapp<=55;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=10729;
 end   
18'd132806: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=5;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=14091;
 end   
18'd132807: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd132808: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd132809: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd132810: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd132811: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd132812: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd132813: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11810;
 end   
18'd132814: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11810;
 end   
18'd132815: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11810;
 end   
18'd132942: begin  
rid<=1;
end
18'd132943: begin  
end
18'd132944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd132945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd132946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd132947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd132948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd132949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd132950: begin  
rid<=0;
end
18'd133001: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=8;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5873;
 end   
18'd133002: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=22;
   mapp<=22;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13777;
 end   
18'd133003: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=40;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd133004: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=1;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd133005: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=37;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd133006: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd133007: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=47;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd133008: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=19;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd133009: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=91;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd133010: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd133011: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd133012: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd133013: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5873;
 end   
18'd133014: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5873;
 end   
18'd133015: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5873;
 end   
18'd133016: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5873;
 end   
18'd133017: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5873;
 end   
18'd133018: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5873;
 end   
18'd133019: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5873;
 end   
18'd133142: begin  
rid<=1;
end
18'd133143: begin  
end
18'd133144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd133145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd133146: begin  
rid<=0;
end
18'd133201: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=25;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=125;
 end   
18'd133202: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=90;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=460;
 end   
18'd133203: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=30;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=170;
 end   
18'd133204: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=81;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=435;
 end   
18'd133205: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=88;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=480;
 end   
18'd133206: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=95;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=525;
 end   
18'd133207: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=38;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=250;
 end   
18'd133208: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd133342: begin  
rid<=1;
end
18'd133343: begin  
end
18'd133344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd133345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd133346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd133347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd133348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd133349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd133350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd133351: begin  
rid<=0;
end
18'd133401: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=1;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12040;
 end   
18'd133402: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=23;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd133403: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=15;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd133404: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=9;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd133405: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=53;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd133406: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=2;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd133407: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=31;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd133408: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=85;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd133409: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=89;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd133410: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd133411: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd133412: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd133413: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12040;
 end   
18'd133414: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12040;
 end   
18'd133415: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12040;
 end   
18'd133416: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12040;
 end   
18'd133417: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12040;
 end   
18'd133418: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12040;
 end   
18'd133542: begin  
rid<=1;
end
18'd133543: begin  
end
18'd133544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd133545: begin  
rid<=0;
end
18'd133601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=38;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11336;
 end   
18'd133602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=55;
   mapp<=64;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10886;
 end   
18'd133603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=15;
   mapp<=12;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=11561;
 end   
18'd133604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=41;
   mapp<=27;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=15597;
 end   
18'd133605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=56;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd133606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=9;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd133607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd133608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd133609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd133610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd133611: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd133612: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd133613: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11336;
 end   
18'd133614: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11336;
 end   
18'd133615: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11336;
 end   
18'd133742: begin  
rid<=1;
end
18'd133743: begin  
end
18'd133744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd133745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd133746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd133747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd133748: begin  
rid<=0;
end
18'd133801: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=31;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12527;
 end   
18'd133802: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=51;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=17418;
 end   
18'd133803: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=51;
   mapp<=79;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=18929;
 end   
18'd133804: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=96;
   mapp<=43;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=18561;
 end   
18'd133805: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=98;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=13168;
 end   
18'd133806: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=79;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=11159;
 end   
18'd133807: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=38;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=9936;
 end   
18'd133808: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=6;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=5448;
 end   
18'd133809: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=91;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd133810: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=1;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd133811: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=13;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd133812: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd133813: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12527;
 end   
18'd133814: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12527;
 end   
18'd133815: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12527;
 end   
18'd133942: begin  
rid<=1;
end
18'd133943: begin  
end
18'd133944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd133945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd133946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd133947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd133948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd133949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd133950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd133951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd133952: begin  
rid<=0;
end
18'd134001: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=35;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=24938;
 end   
18'd134002: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=58;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd134003: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=99;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd134004: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=61;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd134005: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=80;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd134006: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=74;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd134007: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd134008: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd134009: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd134010: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd134011: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd134012: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd134142: begin  
rid<=1;
end
18'd134143: begin  
end
18'd134144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd134145: begin  
rid<=0;
end
18'd134201: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=53;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8372;
 end   
18'd134202: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=99;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13864;
 end   
18'd134203: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=23;
   mapp<=93;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=13809;
 end   
18'd134204: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=73;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=11641;
 end   
18'd134205: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=71;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=8068;
 end   
18'd134206: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd134207: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd134208: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd134209: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd134210: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd134342: begin  
rid<=1;
end
18'd134343: begin  
end
18'd134344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd134345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd134346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd134347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd134348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd134349: begin  
rid<=0;
end
18'd134401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=9;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13796;
 end   
18'd134402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=33;
   mapp<=66;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13569;
 end   
18'd134403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=22;
   mapp<=92;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=13413;
 end   
18'd134404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=82;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd134405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=89;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd134406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=42;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd134407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd134408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd134409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd134410: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd134411: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd134412: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd134413: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13796;
 end   
18'd134414: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13796;
 end   
18'd134542: begin  
rid<=1;
end
18'd134543: begin  
end
18'd134544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd134545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd134546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd134547: begin  
rid<=0;
end
18'd134601: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=65;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2600;
 end   
18'd134602: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=0;
   mapp<=36;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=2350;
 end   
18'd134603: begin  
  clrr<=0;
  maplen<=2;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd134742: begin  
rid<=1;
end
18'd134743: begin  
end
18'd134744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd134745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd134746: begin  
rid<=0;
end
18'd134801: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=96;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=24698;
 end   
18'd134802: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=26;
   mapp<=26;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=22059;
 end   
18'd134803: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=65;
   mapp<=55;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=24862;
 end   
18'd134804: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=85;
   mapp<=25;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=21436;
 end   
18'd134805: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=81;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd134806: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=29;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd134807: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=56;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd134808: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=88;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd134809: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd134810: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd134811: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd134812: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd134813: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24698;
 end   
18'd134814: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24698;
 end   
18'd134815: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24698;
 end   
18'd134816: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24698;
 end   
18'd134817: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24698;
 end   
18'd134818: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24698;
 end   
18'd134819: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24698;
 end   
18'd134942: begin  
rid<=1;
end
18'd134943: begin  
end
18'd134944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd134945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd134946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd134947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd134948: begin  
rid<=0;
end
18'd135001: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=15;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1470;
 end   
18'd135002: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=99;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9712;
 end   
18'd135003: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=22;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=2176;
 end   
18'd135004: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd135142: begin  
rid<=1;
end
18'd135143: begin  
end
18'd135144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd135145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd135146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd135147: begin  
rid<=0;
end
18'd135201: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=16;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1668;
 end   
18'd135202: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=28;
   mapp<=43;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3445;
 end   
18'd135203: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=61;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5659;
 end   
18'd135204: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=90;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=3672;
 end   
18'd135205: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=24;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=2499;
 end   
18'd135206: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=41;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=3260;
 end   
18'd135207: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=47;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=3444;
 end   
18'd135208: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=47;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=2250;
 end   
18'd135209: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=19;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd135210: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd135211: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd135342: begin  
rid<=1;
end
18'd135343: begin  
end
18'd135344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd135345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd135346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd135347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd135348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd135349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd135350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd135351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd135352: begin  
rid<=0;
end
18'd135401: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=68;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=20933;
 end   
18'd135402: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=45;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=17276;
 end   
18'd135403: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=17;
   mapp<=3;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=16635;
 end   
18'd135404: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=45;
   mapp<=49;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=16457;
 end   
18'd135405: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=67;
   mapp<=90;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=13113;
 end   
18'd135406: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=70;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd135407: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd135408: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=86;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd135409: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=25;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd135410: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=2;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd135411: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd135412: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd135413: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20933;
 end   
18'd135414: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20933;
 end   
18'd135415: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20933;
 end   
18'd135416: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20933;
 end   
18'd135542: begin  
rid<=1;
end
18'd135543: begin  
end
18'd135544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd135545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd135546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd135547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd135548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd135549: begin  
rid<=0;
end
18'd135601: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=96;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3788;
 end   
18'd135602: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=20;
   mapp<=55;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2825;
 end   
18'd135603: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=41;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1883;
 end   
18'd135604: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=13;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=2924;
 end   
18'd135605: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=46;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=5618;
 end   
18'd135606: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=78;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=3719;
 end   
18'd135607: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=27;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=981;
 end   
18'd135608: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=3;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=1474;
 end   
18'd135609: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=24;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=5482;
 end   
18'd135610: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=86;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd135611: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd135612: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd135742: begin  
rid<=1;
end
18'd135743: begin  
end
18'd135744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd135745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd135746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd135747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd135748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd135749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd135750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd135751: begin  
check<=expctdoutput[7]-outcheck;
end
18'd135752: begin  
check<=expctdoutput[8]-outcheck;
end
18'd135753: begin  
rid<=0;
end
18'd135801: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=44;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4268;
 end   
18'd135802: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=3002;
 end   
18'd135803: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=16;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=724;
 end   
18'd135804: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=18;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=822;
 end   
18'd135805: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd135942: begin  
rid<=1;
end
18'd135943: begin  
end
18'd135944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd135945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd135946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd135947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd135948: begin  
rid<=0;
end
18'd136001: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=72;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6333;
 end   
18'd136002: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=43;
   mapp<=15;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3512;
 end   
18'd136003: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=7;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=828;
 end   
18'd136004: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=17;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=1763;
 end   
18'd136005: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=26;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=2349;
 end   
18'd136006: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=17;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=2593;
 end   
18'd136007: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=80;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=7235;
 end   
18'd136008: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=57;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd136009: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd136010: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd136142: begin  
rid<=1;
end
18'd136143: begin  
end
18'd136144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd136145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd136146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd136147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd136148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd136149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd136150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd136151: begin  
rid<=0;
end
18'd136201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=35;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6630;
 end   
18'd136202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=28;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10236;
 end   
18'd136203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=14;
   mapp<=22;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5008;
 end   
18'd136204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=58;
   mapp<=74;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=10796;
 end   
18'd136205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=99;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=9360;
 end   
18'd136206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=27;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=5038;
 end   
18'd136207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=92;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd136208: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=21;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd136209: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=40;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd136210: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd136211: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd136212: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd136213: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6630;
 end   
18'd136342: begin  
rid<=1;
end
18'd136343: begin  
end
18'd136344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd136345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd136346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd136347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd136348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd136349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd136350: begin  
rid<=0;
end
18'd136401: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=2;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9544;
 end   
18'd136402: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=43;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6544;
 end   
18'd136403: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=96;
   mapp<=46;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6547;
 end   
18'd136404: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=27;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd136405: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=17;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd136406: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd136407: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd136408: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd136409: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd136410: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd136411: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd136412: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd136542: begin  
rid<=1;
end
18'd136543: begin  
end
18'd136544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd136545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd136546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd136547: begin  
rid<=0;
end
18'd136601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9410;
 end   
18'd136602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=50;
   mapp<=76;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4986;
 end   
18'd136603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=66;
   mapp<=85;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=4926;
 end   
18'd136604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=11;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=6894;
 end   
18'd136605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=66;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=6304;
 end   
18'd136606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=54;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=5522;
 end   
18'd136607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=54;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=4998;
 end   
18'd136608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd136609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd136610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd136611: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd136612: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd136742: begin  
rid<=1;
end
18'd136743: begin  
end
18'd136744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd136745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd136746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd136747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd136748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd136749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd136750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd136751: begin  
rid<=0;
end
18'd136801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=24;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12839;
 end   
18'd136802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=21;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10410;
 end   
18'd136803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=48;
   mapp<=82;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=11402;
 end   
18'd136804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=11;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd136805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=75;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd136806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd136807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd136808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd136809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd136810: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd136811: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd136812: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd136942: begin  
rid<=1;
end
18'd136943: begin  
end
18'd136944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd136945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd136946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd136947: begin  
rid<=0;
end
18'd137001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=4;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=25216;
 end   
18'd137002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=84;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd137003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=81;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd137004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=65;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd137005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=72;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd137006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=30;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd137007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=60;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd137008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=87;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd137009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=15;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd137010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=45;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd137011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=93;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd137012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd137013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25216;
 end   
18'd137014: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25216;
 end   
18'd137015: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25216;
 end   
18'd137016: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25216;
 end   
18'd137017: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25216;
 end   
18'd137018: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25216;
 end   
18'd137019: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25216;
 end   
18'd137020: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25216;
 end   
18'd137021: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25216;
 end   
18'd137022: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25216;
 end   
18'd137142: begin  
rid<=1;
end
18'd137143: begin  
end
18'd137144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd137145: begin  
rid<=0;
end
18'd137201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=66;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13288;
 end   
18'd137202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=70;
   mapp<=49;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11912;
 end   
18'd137203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=96;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd137204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd137205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd137206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd137207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd137342: begin  
rid<=1;
end
18'd137343: begin  
end
18'd137344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd137345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd137346: begin  
rid<=0;
end
18'd137401: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=14;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6940;
 end   
18'd137402: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=24;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4566;
 end   
18'd137403: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=61;
   mapp<=60;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=4255;
 end   
18'd137404: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=25;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd137405: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd137406: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd137407: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd137408: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd137409: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd137410: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd137542: begin  
rid<=1;
end
18'd137543: begin  
end
18'd137544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd137545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd137546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd137547: begin  
rid<=0;
end
18'd137601: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=24;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14111;
 end   
18'd137602: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=46;
   mapp<=49;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=16880;
 end   
18'd137603: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=87;
   mapp<=17;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=18190;
 end   
18'd137604: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=17;
   mapp<=18;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=22213;
 end   
18'd137605: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=82;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd137606: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=71;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd137607: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=40;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd137608: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd137609: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd137610: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd137611: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd137612: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd137613: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14111;
 end   
18'd137614: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14111;
 end   
18'd137615: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14111;
 end   
18'd137616: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14111;
 end   
18'd137617: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14111;
 end   
18'd137742: begin  
rid<=1;
end
18'd137743: begin  
end
18'd137744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd137745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd137746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd137747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd137748: begin  
rid<=0;
end
18'd137801: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=73;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1825;
 end   
18'd137802: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=47;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1185;
 end   
18'd137803: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=6;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=170;
 end   
18'd137804: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=88;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=2230;
 end   
18'd137805: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=17;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=465;
 end   
18'd137806: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=43;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=1125;
 end   
18'd137807: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=38;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=1010;
 end   
18'd137808: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=84;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=2170;
 end   
18'd137809: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=57;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=1505;
 end   
18'd137810: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=39;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[9]<=1065;
 end   
18'd137811: begin  
  clrr<=0;
  maplen<=1;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd137942: begin  
rid<=1;
end
18'd137943: begin  
end
18'd137944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd137945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd137946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd137947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd137948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd137949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd137950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd137951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd137952: begin  
check<=expctdoutput[8]-outcheck;
end
18'd137953: begin  
check<=expctdoutput[9]-outcheck;
end
18'd137954: begin  
rid<=0;
end
18'd138001: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=84;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2604;
 end   
18'd138002: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=53;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=4462;
 end   
18'd138003: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=65;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=5480;
 end   
18'd138004: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=37;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=3138;
 end   
18'd138005: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=90;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=7600;
 end   
18'd138006: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=71;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=6014;
 end   
18'd138007: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=27;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=2328;
 end   
18'd138008: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=97;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=8218;
 end   
18'd138009: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=60;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=5120;
 end   
18'd138010: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd138142: begin  
rid<=1;
end
18'd138143: begin  
end
18'd138144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd138145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd138146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd138147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd138148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd138149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd138150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd138151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd138152: begin  
check<=expctdoutput[8]-outcheck;
end
18'd138153: begin  
rid<=0;
end
18'd138201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=6;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9886;
 end   
18'd138202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=13;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7183;
 end   
18'd138203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=98;
   mapp<=90;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=17958;
 end   
18'd138204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=23;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=11303;
 end   
18'd138205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=90;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=12960;
 end   
18'd138206: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd138207: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=25;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd138208: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd138209: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd138210: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd138342: begin  
rid<=1;
end
18'd138343: begin  
end
18'd138344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd138345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd138346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd138347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd138348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd138349: begin  
rid<=0;
end
18'd138401: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=78;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3588;
 end   
18'd138402: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=78;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=6094;
 end   
18'd138403: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=54;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=4232;
 end   
18'd138404: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=1;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=108;
 end   
18'd138405: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=23;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=1834;
 end   
18'd138406: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=13;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=1064;
 end   
18'd138407: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=98;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=7704;
 end   
18'd138408: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=46;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=3658;
 end   
18'd138409: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=87;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=6866;
 end   
18'd138410: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd138542: begin  
rid<=1;
end
18'd138543: begin  
end
18'd138544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd138545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd138546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd138547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd138548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd138549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd138550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd138551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd138552: begin  
check<=expctdoutput[8]-outcheck;
end
18'd138553: begin  
rid<=0;
end
18'd138601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=26;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16866;
 end   
18'd138602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=92;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd138603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=66;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd138604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=24;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd138605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=44;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd138606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=55;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd138607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=2;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd138608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=19;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd138609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=88;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd138610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd138611: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd138612: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd138613: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16866;
 end   
18'd138614: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16866;
 end   
18'd138615: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16866;
 end   
18'd138616: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16866;
 end   
18'd138617: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16866;
 end   
18'd138618: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16866;
 end   
18'd138742: begin  
rid<=1;
end
18'd138743: begin  
end
18'd138744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd138745: begin  
rid<=0;
end
18'd138801: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=54;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=17904;
 end   
18'd138802: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=2;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=12781;
 end   
18'd138803: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=34;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd138804: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=15;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd138805: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=10;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd138806: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=63;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd138807: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=74;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd138808: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=92;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd138809: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=84;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd138810: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=81;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd138811: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=48;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd138812: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd138813: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17904;
 end   
18'd138814: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17904;
 end   
18'd138815: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17904;
 end   
18'd138816: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17904;
 end   
18'd138817: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17904;
 end   
18'd138818: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17904;
 end   
18'd138819: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17904;
 end   
18'd138820: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17904;
 end   
18'd138821: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17904;
 end   
18'd138942: begin  
rid<=1;
end
18'd138943: begin  
end
18'd138944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd138945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd138946: begin  
rid<=0;
end
18'd139001: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=55;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10143;
 end   
18'd139002: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=79;
   mapp<=81;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=16140;
 end   
18'd139003: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=78;
   mapp<=2;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=18927;
 end   
18'd139004: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=14;
   mapp<=93;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=17745;
 end   
18'd139005: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=7;
   mapp<=96;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=20548;
 end   
18'd139006: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=73;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd139007: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=99;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd139008: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=66;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd139009: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=68;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd139010: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=85;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd139011: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=24;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd139012: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd139013: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10143;
 end   
18'd139014: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10143;
 end   
18'd139015: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10143;
 end   
18'd139016: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10143;
 end   
18'd139017: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10143;
 end   
18'd139018: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10143;
 end   
18'd139142: begin  
rid<=1;
end
18'd139143: begin  
end
18'd139144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd139145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd139146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd139147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd139148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd139149: begin  
rid<=0;
end
18'd139201: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=42;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4076;
 end   
18'd139202: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=97;
   mapp<=18;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3593;
 end   
18'd139203: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=88;
   mapp<=11;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5636;
 end   
18'd139204: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=72;
   mapp<=2;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=12208;
 end   
18'd139205: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd139206: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd139207: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd139208: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd139209: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd139210: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd139211: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd139342: begin  
rid<=1;
end
18'd139343: begin  
end
18'd139344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd139345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd139346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd139347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd139348: begin  
rid<=0;
end
18'd139401: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=9;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1689;
 end   
18'd139402: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=29;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1341;
 end   
18'd139403: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=31;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=1749;
 end   
18'd139404: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=50;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=3264;
 end   
18'd139405: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=96;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=2615;
 end   
18'd139406: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd139407: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd139408: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd139542: begin  
rid<=1;
end
18'd139543: begin  
end
18'd139544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd139545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd139546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd139547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd139548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd139549: begin  
rid<=0;
end
18'd139601: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=38;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=417;
 end   
18'd139602: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=9;
   mapp<=21;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1609;
 end   
18'd139603: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=89;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=3627;
 end   
18'd139604: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd139605: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd139606: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd139742: begin  
rid<=1;
end
18'd139743: begin  
end
18'd139744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd139745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd139746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd139747: begin  
rid<=0;
end
18'd139801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=50;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6032;
 end   
18'd139802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=93;
   mapp<=7;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10054;
 end   
18'd139803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=49;
   mapp<=29;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6882;
 end   
18'd139804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=94;
   mapp<=13;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=11962;
 end   
18'd139805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=2;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd139806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=8;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd139807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd139808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=27;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd139809: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=72;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd139810: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd139811: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd139812: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd139813: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6032;
 end   
18'd139814: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6032;
 end   
18'd139815: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6032;
 end   
18'd139942: begin  
rid<=1;
end
18'd139943: begin  
end
18'd139944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd139945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd139946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd139947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd139948: begin  
rid<=0;
end
18'd140001: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=44;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9774;
 end   
18'd140002: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=58;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6678;
 end   
18'd140003: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=75;
   mapp<=50;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=4109;
 end   
18'd140004: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=8;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=3059;
 end   
18'd140005: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=19;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=8319;
 end   
18'd140006: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=21;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=7813;
 end   
18'd140007: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=83;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=10753;
 end   
18'd140008: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=27;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=5867;
 end   
18'd140009: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd140010: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd140011: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd140012: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd140013: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9774;
 end   
18'd140142: begin  
rid<=1;
end
18'd140143: begin  
end
18'd140144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd140145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd140146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd140147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd140148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd140149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd140150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd140151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd140152: begin  
rid<=0;
end
18'd140201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=86;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8797;
 end   
18'd140202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=63;
   mapp<=52;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5119;
 end   
18'd140203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=31;
   mapp<=83;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6845;
 end   
18'd140204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=1;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd140205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=53;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd140206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=55;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd140207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd140208: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd140209: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd140210: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd140342: begin  
rid<=1;
end
18'd140343: begin  
end
18'd140344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd140345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd140346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd140347: begin  
rid<=0;
end
18'd140401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=91;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6009;
 end   
18'd140402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=52;
   mapp<=51;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9993;
 end   
18'd140403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=9;
   mapp<=61;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8189;
 end   
18'd140404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=26;
   mapp<=10;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=6279;
 end   
18'd140405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=80;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=12685;
 end   
18'd140406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd140407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd140408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd140409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd140410: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd140411: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd140412: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd140542: begin  
rid<=1;
end
18'd140543: begin  
end
18'd140544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd140545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd140546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd140547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd140548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd140549: begin  
rid<=0;
end
18'd140601: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=21;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3333;
 end   
18'd140602: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=67;
   mapp<=30;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5701;
 end   
18'd140603: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=49;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=3617;
 end   
18'd140604: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=17;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=3051;
 end   
18'd140605: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=65;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=4465;
 end   
18'd140606: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=11;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=1493;
 end   
18'd140607: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=25;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=1875;
 end   
18'd140608: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=8;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=2434;
 end   
18'd140609: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd140610: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd140611: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd140742: begin  
rid<=1;
end
18'd140743: begin  
end
18'd140744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd140745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd140746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd140747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd140748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd140749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd140750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd140751: begin  
check<=expctdoutput[7]-outcheck;
end
18'd140752: begin  
rid<=0;
end
18'd140801: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=21;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14697;
 end   
18'd140802: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=80;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd140803: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=37;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd140804: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=69;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd140805: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=7;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd140806: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd140807: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd140808: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd140809: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd140810: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd140942: begin  
rid<=1;
end
18'd140943: begin  
end
18'd140944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd140945: begin  
rid<=0;
end
18'd141001: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=70;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=24157;
 end   
18'd141002: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=59;
   mapp<=82;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=20339;
 end   
18'd141003: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=33;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd141004: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=56;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd141005: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=93;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd141006: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=91;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd141007: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd141008: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd141009: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd141010: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd141011: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd141012: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd141013: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24157;
 end   
18'd141142: begin  
rid<=1;
end
18'd141143: begin  
end
18'd141144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd141145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd141146: begin  
rid<=0;
end
18'd141201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=28;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7018;
 end   
18'd141202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=46;
   mapp<=57;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=14658;
 end   
18'd141203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=20;
   mapp<=98;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=10131;
 end   
18'd141204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=97;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=17374;
 end   
18'd141205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=29;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=15503;
 end   
18'd141206: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=74;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=17343;
 end   
18'd141207: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=89;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=17438;
 end   
18'd141208: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=59;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd141209: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=64;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd141210: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd141211: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd141212: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd141342: begin  
rid<=1;
end
18'd141343: begin  
end
18'd141344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd141345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd141346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd141347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd141348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd141349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd141350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd141351: begin  
rid<=0;
end
18'd141401: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=78;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12519;
 end   
18'd141402: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=54;
   mapp<=8;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10666;
 end   
18'd141403: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=64;
   mapp<=17;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9619;
 end   
18'd141404: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=47;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd141405: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=3;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd141406: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=24;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd141407: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=26;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd141408: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd141409: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd141410: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd141411: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd141412: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd141413: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12519;
 end   
18'd141414: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12519;
 end   
18'd141415: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12519;
 end   
18'd141416: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12519;
 end   
18'd141542: begin  
rid<=1;
end
18'd141543: begin  
end
18'd141544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd141545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd141546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd141547: begin  
rid<=0;
end
18'd141601: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=75;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9200;
 end   
18'd141602: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=25;
   mapp<=92;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8260;
 end   
18'd141603: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=54;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=4820;
 end   
18'd141604: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=30;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=3505;
 end   
18'd141605: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd141606: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd141607: begin  
  clrr<=0;
  maplen<=5;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd141742: begin  
rid<=1;
end
18'd141743: begin  
end
18'd141744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd141745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd141746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd141747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd141748: begin  
rid<=0;
end
18'd141801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=37;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5134;
 end   
18'd141802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=40;
   mapp<=71;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8738;
 end   
18'd141803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=88;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9310;
 end   
18'd141804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=54;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=7851;
 end   
18'd141805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=63;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=8703;
 end   
18'd141806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=67;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd141807: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd141808: begin  
  clrr<=0;
  maplen<=2;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd141942: begin  
rid<=1;
end
18'd141943: begin  
end
18'd141944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd141945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd141946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd141947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd141948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd141949: begin  
rid<=0;
end
18'd142001: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=72;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8956;
 end   
18'd142002: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=53;
   mapp<=13;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8010;
 end   
18'd142003: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=65;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd142004: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=45;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd142005: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=6;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd142006: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=26;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd142007: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=57;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd142008: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=96;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd142009: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd142010: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd142011: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd142012: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd142013: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8956;
 end   
18'd142014: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8956;
 end   
18'd142015: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8956;
 end   
18'd142142: begin  
rid<=1;
end
18'd142143: begin  
end
18'd142144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd142145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd142146: begin  
rid<=0;
end
18'd142201: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=56;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=20940;
 end   
18'd142202: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=79;
   mapp<=84;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=21085;
 end   
18'd142203: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=96;
   mapp<=93;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=13134;
 end   
18'd142204: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=94;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=11353;
 end   
18'd142205: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=5;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=8629;
 end   
18'd142206: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd142207: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd142208: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd142209: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd142210: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd142342: begin  
rid<=1;
end
18'd142343: begin  
end
18'd142344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd142345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd142346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd142347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd142348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd142349: begin  
rid<=0;
end
18'd142401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=36;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5334;
 end   
18'd142402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=79;
   mapp<=42;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4682;
 end   
18'd142403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd142404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd142405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd142542: begin  
rid<=1;
end
18'd142543: begin  
end
18'd142544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd142545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd142546: begin  
rid<=0;
end
18'd142601: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=32;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=192;
 end   
18'd142602: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=79;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=484;
 end   
18'd142603: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=90;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=560;
 end   
18'd142604: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=35;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=240;
 end   
18'd142605: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd142742: begin  
rid<=1;
end
18'd142743: begin  
end
18'd142744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd142745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd142746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd142747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd142748: begin  
rid<=0;
end
18'd142801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=17;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7003;
 end   
18'd142802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=78;
   mapp<=73;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6235;
 end   
18'd142803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=3;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6164;
 end   
18'd142804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=81;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd142805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd142806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd142942: begin  
rid<=1;
end
18'd142943: begin  
end
18'd142944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd142945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd142946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd142947: begin  
rid<=0;
end
18'd143001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=61;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13088;
 end   
18'd143002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=97;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=12232;
 end   
18'd143003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=53;
   mapp<=40;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9516;
 end   
18'd143004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=9;
   mapp<=31;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=7510;
 end   
18'd143005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=35;
   mapp<=86;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=8988;
 end   
18'd143006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=21;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=6068;
 end   
18'd143007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd143008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=43;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd143009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=33;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd143010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=6;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd143011: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd143012: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd143013: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13088;
 end   
18'd143014: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13088;
 end   
18'd143015: begin  
  clrr<=0;
  maplen<=5;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13088;
 end   
18'd143142: begin  
rid<=1;
end
18'd143143: begin  
end
18'd143144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd143145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd143146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd143147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd143148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd143149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd143150: begin  
rid<=0;
end
18'd143201: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=52;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5504;
 end   
18'd143202: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=26;
   mapp<=73;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5926;
 end   
18'd143203: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=31;
   mapp<=34;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6804;
 end   
18'd143204: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=69;
   mapp<=7;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=4650;
 end   
18'd143205: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=8;
   mapp<=4;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=4416;
 end   
18'd143206: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=31;
   mapp<=7;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=4564;
 end   
18'd143207: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=31;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd143208: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=7;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd143209: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=46;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd143210: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=78;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd143211: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=42;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd143212: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd143213: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5504;
 end   
18'd143214: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5504;
 end   
18'd143215: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5504;
 end   
18'd143216: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5504;
 end   
18'd143217: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5504;
 end   
18'd143342: begin  
rid<=1;
end
18'd143343: begin  
end
18'd143344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd143345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd143346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd143347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd143348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd143349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd143350: begin  
rid<=0;
end
18'd143401: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=14;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11915;
 end   
18'd143402: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=86;
   mapp<=47;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11738;
 end   
18'd143403: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=5;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd143404: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=39;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd143405: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=65;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd143406: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=21;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd143407: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd143408: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd143409: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd143410: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd143411: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd143542: begin  
rid<=1;
end
18'd143543: begin  
end
18'd143544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd143545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd143546: begin  
rid<=0;
end
18'd143601: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=16;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1672;
 end   
18'd143602: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=38;
   mapp<=20;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2796;
 end   
18'd143603: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=31;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=3547;
 end   
18'd143604: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=88;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=5926;
 end   
18'd143605: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=44;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd143606: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd143607: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd143742: begin  
rid<=1;
end
18'd143743: begin  
end
18'd143744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd143745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd143746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd143747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd143748: begin  
rid<=0;
end
18'd143801: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=88;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=88;
 end   
18'd143802: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd143942: begin  
rid<=1;
end
18'd143943: begin  
end
18'd143944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd143945: begin  
rid<=0;
end
18'd144001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=5;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8578;
 end   
18'd144002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=30;
   mapp<=34;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13140;
 end   
18'd144003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=31;
   mapp<=41;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8557;
 end   
18'd144004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=10;
   mapp<=65;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=6065;
 end   
18'd144005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=5;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd144006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=97;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd144007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=18;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd144008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=16;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd144009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd144010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd144011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd144012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd144013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8578;
 end   
18'd144014: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8578;
 end   
18'd144015: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8578;
 end   
18'd144016: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8578;
 end   
18'd144017: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8578;
 end   
18'd144018: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8578;
 end   
18'd144019: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8578;
 end   
18'd144142: begin  
rid<=1;
end
18'd144143: begin  
end
18'd144144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd144145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd144146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd144147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd144148: begin  
rid<=0;
end
18'd144201: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=18;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=594;
 end   
18'd144202: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=3;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=109;
 end   
18'd144203: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=11;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=383;
 end   
18'd144204: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=60;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=2010;
 end   
18'd144205: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=35;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=1195;
 end   
18'd144206: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=90;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=3020;
 end   
18'd144207: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=20;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=720;
 end   
18'd144208: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd144342: begin  
rid<=1;
end
18'd144343: begin  
end
18'd144344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd144345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd144346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd144347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd144348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd144349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd144350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd144351: begin  
rid<=0;
end
18'd144401: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=68;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10692;
 end   
18'd144402: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=6;
   mapp<=90;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8444;
 end   
18'd144403: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=7;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd144404: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=56;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd144405: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=1;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd144406: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=79;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd144407: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd144408: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd144409: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd144410: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd144411: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd144412: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd144413: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10692;
 end   
18'd144542: begin  
rid<=1;
end
18'd144543: begin  
end
18'd144544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd144545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd144546: begin  
rid<=0;
end
18'd144601: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=33;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3902;
 end   
18'd144602: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=48;
   mapp<=13;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4923;
 end   
18'd144603: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=30;
   mapp<=46;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9476;
 end   
18'd144604: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=4;
   mapp<=43;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=8499;
 end   
18'd144605: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=62;
   mapp<=14;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=10206;
 end   
18'd144606: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=15;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=12087;
 end   
18'd144607: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd144608: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd144609: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd144610: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd144611: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd144612: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd144613: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=3902;
 end   
18'd144614: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=3902;
 end   
18'd144615: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=3902;
 end   
18'd144742: begin  
rid<=1;
end
18'd144743: begin  
end
18'd144744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd144745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd144746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd144747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd144748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd144749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd144750: begin  
rid<=0;
end
18'd144801: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=68;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2712;
 end   
18'd144802: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=30;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd144803: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=38;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd144804: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd144805: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd144806: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd144942: begin  
rid<=1;
end
18'd144943: begin  
end
18'd144944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd144945: begin  
rid<=0;
end
18'd145001: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=65;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8430;
 end   
18'd145002: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=37;
   mapp<=91;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11342;
 end   
18'd145003: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=19;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd145004: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=18;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd145005: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=49;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd145006: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=12;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd145007: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd145008: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd145009: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd145010: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd145011: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd145012: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd145013: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8430;
 end   
18'd145142: begin  
rid<=1;
end
18'd145143: begin  
end
18'd145144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd145145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd145146: begin  
rid<=0;
end
18'd145201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=33;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15672;
 end   
18'd145202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=72;
   mapp<=89;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=15437;
 end   
18'd145203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=89;
   mapp<=90;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12079;
 end   
18'd145204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=53;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=11810;
 end   
18'd145205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=44;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=7767;
 end   
18'd145206: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=65;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=9087;
 end   
18'd145207: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=3;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=12614;
 end   
18'd145208: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=70;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd145209: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=69;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd145210: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd145211: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd145212: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd145342: begin  
rid<=1;
end
18'd145343: begin  
end
18'd145344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd145345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd145346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd145347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd145348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd145349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd145350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd145351: begin  
rid<=0;
end
18'd145401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=88;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10216;
 end   
18'd145402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=66;
   mapp<=24;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8004;
 end   
18'd145403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=96;
   mapp<=56;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9780;
 end   
18'd145404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=58;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd145405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=86;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd145406: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd145407: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd145408: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd145542: begin  
rid<=1;
end
18'd145543: begin  
end
18'd145544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd145545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd145546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd145547: begin  
rid<=0;
end
18'd145601: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=21;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=18803;
 end   
18'd145602: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=87;
   mapp<=76;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=12105;
 end   
18'd145603: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=9;
   mapp<=9;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=13321;
 end   
18'd145604: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=89;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd145605: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=83;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd145606: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=21;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd145607: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=87;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd145608: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd145609: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd145610: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd145611: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd145612: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd145742: begin  
rid<=1;
end
18'd145743: begin  
end
18'd145744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd145745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd145746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd145747: begin  
rid<=0;
end
18'd145801: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=14;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=532;
 end   
18'd145802: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=62;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2366;
 end   
18'd145803: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=55;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=2110;
 end   
18'd145804: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=77;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=2956;
 end   
18'd145805: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=6;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=268;
 end   
18'd145806: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=19;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=772;
 end   
18'd145807: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=43;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=1694;
 end   
18'd145808: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=2;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=146;
 end   
18'd145809: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=12;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=536;
 end   
18'd145810: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=21;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[9]<=888;
 end   
18'd145811: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=92;
   mapp<=0;
   pp<=100;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[10]<=3596;
 end   
18'd145812: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd145942: begin  
rid<=1;
end
18'd145943: begin  
end
18'd145944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd145945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd145946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd145947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd145948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd145949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd145950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd145951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd145952: begin  
check<=expctdoutput[8]-outcheck;
end
18'd145953: begin  
check<=expctdoutput[9]-outcheck;
end
18'd145954: begin  
check<=expctdoutput[10]-outcheck;
end
18'd145955: begin  
rid<=0;
end
18'd146001: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=48;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2112;
 end   
18'd146002: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=15;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=670;
 end   
18'd146003: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=79;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=3496;
 end   
18'd146004: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=21;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=954;
 end   
18'd146005: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=48;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=2152;
 end   
18'd146006: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=51;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=2294;
 end   
18'd146007: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=87;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=3888;
 end   
18'd146008: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=75;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=3370;
 end   
18'd146009: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=79;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=3556;
 end   
18'd146010: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd146142: begin  
rid<=1;
end
18'd146143: begin  
end
18'd146144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd146145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd146146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd146147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd146148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd146149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd146150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd146151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd146152: begin  
check<=expctdoutput[8]-outcheck;
end
18'd146153: begin  
rid<=0;
end
18'd146201: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=87;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4002;
 end   
18'd146202: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=7;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=332;
 end   
18'd146203: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=88;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=4068;
 end   
18'd146204: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=25;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=1180;
 end   
18'd146205: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=95;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=4410;
 end   
18'd146206: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd146342: begin  
rid<=1;
end
18'd146343: begin  
end
18'd146344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd146345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd146346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd146347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd146348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd146349: begin  
rid<=0;
end
18'd146401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=54;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12260;
 end   
18'd146402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=72;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=12708;
 end   
18'd146403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=46;
   mapp<=56;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12336;
 end   
18'd146404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=56;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=10363;
 end   
18'd146405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=79;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=12358;
 end   
18'd146406: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=6449;
 end   
18'd146407: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=93;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=9135;
 end   
18'd146408: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=3;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=1391;
 end   
18'd146409: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=9;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=6186;
 end   
18'd146410: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=8;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd146411: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=85;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd146412: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd146413: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12260;
 end   
18'd146414: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12260;
 end   
18'd146542: begin  
rid<=1;
end
18'd146543: begin  
end
18'd146544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd146545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd146546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd146547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd146548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd146549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd146550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd146551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd146552: begin  
check<=expctdoutput[8]-outcheck;
end
18'd146553: begin  
rid<=0;
end
18'd146601: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=50;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5107;
 end   
18'd146602: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=41;
   mapp<=27;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3344;
 end   
18'd146603: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=2;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=2691;
 end   
18'd146604: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=93;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd146605: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd146606: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd146742: begin  
rid<=1;
end
18'd146743: begin  
end
18'd146744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd146745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd146746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd146747: begin  
rid<=0;
end
18'd146801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=3;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3759;
 end   
18'd146802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=66;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2964;
 end   
18'd146803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=28;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5536;
 end   
18'd146804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=88;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=2550;
 end   
18'd146805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=12;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=3876;
 end   
18'd146806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=64;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=3354;
 end   
18'd146807: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=35;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=4827;
 end   
18'd146808: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=72;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=3430;
 end   
18'd146809: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=33;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=1893;
 end   
18'd146810: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=20;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd146811: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd146812: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd146942: begin  
rid<=1;
end
18'd146943: begin  
end
18'd146944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd146945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd146946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd146947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd146948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd146949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd146950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd146951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd146952: begin  
check<=expctdoutput[8]-outcheck;
end
18'd146953: begin  
rid<=0;
end
18'd147001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=84;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10772;
 end   
18'd147002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=64;
   mapp<=6;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10247;
 end   
18'd147003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=85;
   mapp<=13;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6834;
 end   
18'd147004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=71;
   mapp<=61;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=7354;
 end   
18'd147005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=92;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd147006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd147007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd147008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd147009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd147010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd147011: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd147012: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd147013: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10772;
 end   
18'd147142: begin  
rid<=1;
end
18'd147143: begin  
end
18'd147144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd147145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd147146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd147147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd147148: begin  
rid<=0;
end
18'd147201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=67;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15343;
 end   
18'd147202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=38;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd147203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=56;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd147204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=98;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd147205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd147206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd147207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd147208: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd147342: begin  
rid<=1;
end
18'd147343: begin  
end
18'd147344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd147345: begin  
rid<=0;
end
18'd147401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=27;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7791;
 end   
18'd147402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=3;
   mapp<=64;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13813;
 end   
18'd147403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=55;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd147404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=39;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd147405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=40;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd147406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=19;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd147407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=80;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd147408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=93;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd147409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=57;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd147410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=92;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd147411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd147412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd147413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7791;
 end   
18'd147414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7791;
 end   
18'd147415: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7791;
 end   
18'd147416: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7791;
 end   
18'd147417: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7791;
 end   
18'd147418: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7791;
 end   
18'd147419: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7791;
 end   
18'd147420: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7791;
 end   
18'd147421: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7791;
 end   
18'd147542: begin  
rid<=1;
end
18'd147543: begin  
end
18'd147544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd147545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd147546: begin  
rid<=0;
end
18'd147601: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=42;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6126;
 end   
18'd147602: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=79;
   mapp<=39;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8411;
 end   
18'd147603: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=7;
   mapp<=81;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8111;
 end   
18'd147604: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd147605: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd147606: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd147607: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd147608: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd147742: begin  
rid<=1;
end
18'd147743: begin  
end
18'd147744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd147745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd147746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd147747: begin  
rid<=0;
end
18'd147801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=94;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11339;
 end   
18'd147802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=63;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5184;
 end   
18'd147803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=13;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=2940;
 end   
18'd147804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=25;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=6718;
 end   
18'd147805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=61;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=12056;
 end   
18'd147806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=97;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=11418;
 end   
18'd147807: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=61;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=11080;
 end   
18'd147808: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=85;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd147809: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd147810: begin  
  clrr<=0;
  maplen<=2;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd147942: begin  
rid<=1;
end
18'd147943: begin  
end
18'd147944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd147945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd147946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd147947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd147948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd147949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd147950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd147951: begin  
rid<=0;
end
18'd148001: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=50;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16192;
 end   
18'd148002: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=85;
   mapp<=44;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=14133;
 end   
18'd148003: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=20;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd148004: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=31;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd148005: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=16;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd148006: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=86;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd148007: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd148008: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd148009: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd148010: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd148011: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd148012: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd148013: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16192;
 end   
18'd148142: begin  
rid<=1;
end
18'd148143: begin  
end
18'd148144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd148145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd148146: begin  
rid<=0;
end
18'd148201: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=47;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=799;
 end   
18'd148202: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=89;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1523;
 end   
18'd148203: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=92;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1584;
 end   
18'd148204: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=96;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=1662;
 end   
18'd148205: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd148342: begin  
rid<=1;
end
18'd148343: begin  
end
18'd148344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd148345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd148346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd148347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd148348: begin  
rid<=0;
end
18'd148401: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=61;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=17612;
 end   
18'd148402: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=81;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=16096;
 end   
18'd148403: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=41;
   mapp<=23;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=17320;
 end   
18'd148404: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=61;
   mapp<=91;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=18171;
 end   
18'd148405: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=43;
   mapp<=66;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=14961;
 end   
18'd148406: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=45;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd148407: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=96;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd148408: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=29;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd148409: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=73;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd148410: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd148411: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd148412: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd148413: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17612;
 end   
18'd148414: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17612;
 end   
18'd148542: begin  
rid<=1;
end
18'd148543: begin  
end
18'd148544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd148545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd148546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd148547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd148548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd148549: begin  
rid<=0;
end
18'd148601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=88;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11588;
 end   
18'd148602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=79;
   mapp<=28;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7852;
 end   
18'd148603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=73;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd148604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=20;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd148605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=37;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd148606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=55;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd148607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=14;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd148608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=31;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd148609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd148610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=97;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd148611: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd148612: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd148613: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11588;
 end   
18'd148614: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11588;
 end   
18'd148615: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11588;
 end   
18'd148616: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11588;
 end   
18'd148617: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11588;
 end   
18'd148618: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11588;
 end   
18'd148619: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11588;
 end   
18'd148742: begin  
rid<=1;
end
18'd148743: begin  
end
18'd148744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd148745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd148746: begin  
rid<=0;
end
18'd148801: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=29;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=603;
 end   
18'd148802: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=13;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=567;
 end   
18'd148803: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=3;
   mapp<=28;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1534;
 end   
18'd148804: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=45;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=1929;
 end   
18'd148805: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=39;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=1845;
 end   
18'd148806: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=29;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=2277;
 end   
18'd148807: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=99;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=3648;
 end   
18'd148808: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=33;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=2527;
 end   
18'd148809: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=96;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=4184;
 end   
18'd148810: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd148811: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd148812: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd148813: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=603;
 end   
18'd148814: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=603;
 end   
18'd148942: begin  
rid<=1;
end
18'd148943: begin  
end
18'd148944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd148945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd148946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd148947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd148948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd148949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd148950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd148951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd148952: begin  
check<=expctdoutput[8]-outcheck;
end
18'd148953: begin  
rid<=0;
end
18'd149001: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=98;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10262;
 end   
18'd149002: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=42;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd149003: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd149004: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd149142: begin  
rid<=1;
end
18'd149143: begin  
end
18'd149144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd149145: begin  
rid<=0;
end
18'd149201: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=70;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14609;
 end   
18'd149202: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=49;
   mapp<=22;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=12713;
 end   
18'd149203: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=97;
   mapp<=15;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=13579;
 end   
18'd149204: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=91;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd149205: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=24;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd149206: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=52;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd149207: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=21;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd149208: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd149209: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd149210: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd149211: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd149212: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd149342: begin  
rid<=1;
end
18'd149343: begin  
end
18'd149344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd149345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd149346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd149347: begin  
rid<=0;
end
18'd149401: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=89;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4651;
 end   
18'd149402: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=96;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd149403: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd149404: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd149542: begin  
rid<=1;
end
18'd149543: begin  
end
18'd149544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd149545: begin  
rid<=0;
end
18'd149601: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=70;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11829;
 end   
18'd149602: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=62;
   mapp<=43;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13082;
 end   
18'd149603: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=63;
   mapp<=81;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=11091;
 end   
18'd149604: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=80;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=8332;
 end   
18'd149605: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd149606: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd149607: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd149608: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd149609: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd149742: begin  
rid<=1;
end
18'd149743: begin  
end
18'd149744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd149745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd149746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd149747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd149748: begin  
rid<=0;
end
18'd149801: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=61;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11322;
 end   
18'd149802: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=98;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13595;
 end   
18'd149803: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=93;
   mapp<=72;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=14045;
 end   
18'd149804: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=41;
   mapp<=31;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=11402;
 end   
18'd149805: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=49;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=12253;
 end   
18'd149806: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=44;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd149807: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd149808: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=82;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd149809: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd149810: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd149811: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd149812: begin  
  clrr<=0;
  maplen<=4;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd149942: begin  
rid<=1;
end
18'd149943: begin  
end
18'd149944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd149945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd149946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd149947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd149948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd149949: begin  
rid<=0;
end
18'd150001: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=6;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6737;
 end   
18'd150002: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=47;
   mapp<=16;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=15576;
 end   
18'd150003: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=6;
   mapp<=10;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=10933;
 end   
18'd150004: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=52;
   mapp<=42;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=10631;
 end   
18'd150005: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=96;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd150006: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=71;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd150007: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd150008: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=77;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd150009: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=56;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd150010: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=35;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd150011: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=11;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd150012: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd150013: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6737;
 end   
18'd150014: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6737;
 end   
18'd150015: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6737;
 end   
18'd150016: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6737;
 end   
18'd150017: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6737;
 end   
18'd150018: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6737;
 end   
18'd150019: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6737;
 end   
18'd150142: begin  
rid<=1;
end
18'd150143: begin  
end
18'd150144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd150145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd150146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd150147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd150148: begin  
rid<=0;
end
18'd150201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=32;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11311;
 end   
18'd150202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=79;
   mapp<=23;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8740;
 end   
18'd150203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=82;
   mapp<=83;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8990;
 end   
18'd150204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=13;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=5771;
 end   
18'd150205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=16;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=6378;
 end   
18'd150206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=58;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=6609;
 end   
18'd150207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=43;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd150208: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=7;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd150209: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=9;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd150210: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd150211: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd150212: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd150213: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11311;
 end   
18'd150342: begin  
rid<=1;
end
18'd150343: begin  
end
18'd150344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd150345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd150346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd150347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd150348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd150349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd150350: begin  
rid<=0;
end
18'd150401: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=7;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13116;
 end   
18'd150402: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=11;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=16652;
 end   
18'd150403: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=57;
   mapp<=17;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=16137;
 end   
18'd150404: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=93;
   mapp<=58;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=14779;
 end   
18'd150405: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=71;
   mapp<=81;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=12789;
 end   
18'd150406: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd150407: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd150408: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd150409: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd150410: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd150411: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd150412: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd150413: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13116;
 end   
18'd150414: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13116;
 end   
18'd150542: begin  
rid<=1;
end
18'd150543: begin  
end
18'd150544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd150545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd150546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd150547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd150548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd150549: begin  
rid<=0;
end
18'd150601: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=77;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=24712;
 end   
18'd150602: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=57;
   mapp<=2;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=20992;
 end   
18'd150603: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=85;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd150604: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=93;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd150605: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=16;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd150606: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=28;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd150607: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=94;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd150608: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd150609: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd150610: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd150611: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd150612: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd150613: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24712;
 end   
18'd150742: begin  
rid<=1;
end
18'd150743: begin  
end
18'd150744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd150745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd150746: begin  
rid<=0;
end
18'd150801: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=91;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9846;
 end   
18'd150802: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=83;
   mapp<=12;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13022;
 end   
18'd150803: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=81;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd150804: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=70;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd150805: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=32;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd150806: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=4;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd150807: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=18;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd150808: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=14;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd150809: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=13;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd150810: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=74;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd150811: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd150812: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd150813: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9846;
 end   
18'd150814: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9846;
 end   
18'd150815: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9846;
 end   
18'd150816: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9846;
 end   
18'd150817: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9846;
 end   
18'd150818: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9846;
 end   
18'd150819: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9846;
 end   
18'd150942: begin  
rid<=1;
end
18'd150943: begin  
end
18'd150944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd150945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd150946: begin  
rid<=0;
end
18'd151001: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=84;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11989;
 end   
18'd151002: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=77;
   mapp<=15;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=12891;
 end   
18'd151003: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=46;
   mapp<=37;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=18496;
 end   
18'd151004: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=20;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd151005: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=6;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd151006: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=62;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd151007: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd151008: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd151009: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd151010: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd151011: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd151012: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd151013: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11989;
 end   
18'd151014: begin  
  clrr<=0;
  maplen<=8;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11989;
 end   
18'd151142: begin  
rid<=1;
end
18'd151143: begin  
end
18'd151144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd151145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd151146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd151147: begin  
rid<=0;
end
18'd151201: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=39;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3231;
 end   
18'd151202: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=51;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4216;
 end   
18'd151203: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=58;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=7076;
 end   
18'd151204: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=94;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=6450;
 end   
18'd151205: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=54;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=6940;
 end   
18'd151206: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=94;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=4379;
 end   
18'd151207: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=13;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=2505;
 end   
18'd151208: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=38;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=6550;
 end   
18'd151209: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=98;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=4157;
 end   
18'd151210: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd151211: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd151212: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd151342: begin  
rid<=1;
end
18'd151343: begin  
end
18'd151344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd151345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd151346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd151347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd151348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd151349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd151350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd151351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd151352: begin  
check<=expctdoutput[8]-outcheck;
end
18'd151353: begin  
rid<=0;
end
18'd151401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=41;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=21441;
 end   
18'd151402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=25;
   mapp<=79;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=26055;
 end   
18'd151403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=40;
   mapp<=17;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=29250;
 end   
18'd151404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=99;
   mapp<=45;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=22619;
 end   
18'd151405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=9;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd151406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=56;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd151407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=43;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd151408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=92;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd151409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=90;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd151410: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=74;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd151411: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=58;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd151412: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd151413: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21441;
 end   
18'd151414: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21441;
 end   
18'd151415: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21441;
 end   
18'd151416: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21441;
 end   
18'd151417: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21441;
 end   
18'd151418: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21441;
 end   
18'd151419: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21441;
 end   
18'd151542: begin  
rid<=1;
end
18'd151543: begin  
end
18'd151544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd151545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd151546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd151547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd151548: begin  
rid<=0;
end
18'd151601: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=0;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=0;
 end   
18'd151602: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=64;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4682;
 end   
18'd151603: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=54;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=3962;
 end   
18'd151604: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=67;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=4921;
 end   
18'd151605: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd151742: begin  
rid<=1;
end
18'd151743: begin  
end
18'd151744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd151745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd151746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd151747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd151748: begin  
rid<=0;
end
18'd151801: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=34;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10429;
 end   
18'd151802: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=20;
   mapp<=75;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9796;
 end   
18'd151803: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=93;
   mapp<=77;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9661;
 end   
18'd151804: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=23;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=8769;
 end   
18'd151805: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=40;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=7931;
 end   
18'd151806: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=59;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=6624;
 end   
18'd151807: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=18;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=8948;
 end   
18'd151808: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=28;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=10691;
 end   
18'd151809: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=76;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd151810: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=45;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd151811: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd151812: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd151813: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10429;
 end   
18'd151942: begin  
rid<=1;
end
18'd151943: begin  
end
18'd151944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd151945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd151946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd151947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd151948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd151949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd151950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd151951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd151952: begin  
rid<=0;
end
18'd152001: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=80;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10726;
 end   
18'd152002: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=26;
   mapp<=26;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8358;
 end   
18'd152003: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=59;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=10805;
 end   
18'd152004: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=60;
   mapp<=12;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=6820;
 end   
18'd152005: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=77;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=11221;
 end   
18'd152006: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=8756;
 end   
18'd152007: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=74;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd152008: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=83;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd152009: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=81;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd152010: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd152011: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd152012: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd152013: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10726;
 end   
18'd152142: begin  
rid<=1;
end
18'd152143: begin  
end
18'd152144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd152145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd152146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd152147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd152148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd152149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd152150: begin  
rid<=0;
end
18'd152201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=41;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9449;
 end   
18'd152202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=5;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9587;
 end   
18'd152203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=94;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd152204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=30;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd152205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=30;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd152206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd152207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd152208: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd152209: begin  
  clrr<=0;
  maplen<=4;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd152342: begin  
rid<=1;
end
18'd152343: begin  
end
18'd152344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd152345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd152346: begin  
rid<=0;
end
18'd152401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=67;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2613;
 end   
18'd152402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=46;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=3092;
 end   
18'd152403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=62;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=4174;
 end   
18'd152404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd152542: begin  
rid<=1;
end
18'd152543: begin  
end
18'd152544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd152545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd152546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd152547: begin  
rid<=0;
end
18'd152601: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=14;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4442;
 end   
18'd152602: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=87;
   mapp<=30;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8038;
 end   
18'd152603: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=60;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd152604: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd152605: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd152606: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd152607: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd152742: begin  
rid<=1;
end
18'd152743: begin  
end
18'd152744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd152745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd152746: begin  
rid<=0;
end
18'd152801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=70;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=20961;
 end   
18'd152802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=55;
   mapp<=43;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=17105;
 end   
18'd152803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=60;
   mapp<=19;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=16490;
 end   
18'd152804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=8;
   mapp<=26;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=12771;
 end   
18'd152805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=98;
   mapp<=48;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=16557;
 end   
18'd152806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=63;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd152807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=84;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd152808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=25;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd152809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=58;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd152810: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=14;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd152811: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=30;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd152812: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd152813: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20961;
 end   
18'd152814: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20961;
 end   
18'd152815: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20961;
 end   
18'd152816: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20961;
 end   
18'd152817: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20961;
 end   
18'd152818: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20961;
 end   
18'd152942: begin  
rid<=1;
end
18'd152943: begin  
end
18'd152944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd152945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd152946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd152947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd152948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd152949: begin  
rid<=0;
end
18'd153001: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=60;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12587;
 end   
18'd153002: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=29;
   mapp<=85;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11731;
 end   
18'd153003: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=43;
   mapp<=0;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=10381;
 end   
18'd153004: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=82;
   mapp<=51;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=15312;
 end   
18'd153005: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=54;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=10040;
 end   
18'd153006: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=80;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=12010;
 end   
18'd153007: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd153008: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd153009: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd153010: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd153011: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd153012: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd153013: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12587;
 end   
18'd153142: begin  
rid<=1;
end
18'd153143: begin  
end
18'd153144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd153145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd153146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd153147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd153148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd153149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd153150: begin  
rid<=0;
end
18'd153201: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=41;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16328;
 end   
18'd153202: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=44;
   mapp<=80;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=20481;
 end   
18'd153203: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=75;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd153204: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=72;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd153205: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=33;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd153206: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=94;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd153207: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd153208: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd153209: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd153210: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd153211: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd153342: begin  
rid<=1;
end
18'd153343: begin  
end
18'd153344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd153345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd153346: begin  
rid<=0;
end
18'd153401: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=77;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12191;
 end   
18'd153402: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=89;
   mapp<=26;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13515;
 end   
18'd153403: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=50;
   mapp<=45;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9782;
 end   
18'd153404: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=78;
   mapp<=4;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=12435;
 end   
18'd153405: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=60;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=10302;
 end   
18'd153406: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=71;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=8599;
 end   
18'd153407: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=60;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=6972;
 end   
18'd153408: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=4;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=5583;
 end   
18'd153409: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd153410: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=97;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd153411: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd153412: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd153413: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12191;
 end   
18'd153414: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12191;
 end   
18'd153415: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12191;
 end   
18'd153542: begin  
rid<=1;
end
18'd153543: begin  
end
18'd153544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd153545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd153546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd153547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd153548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd153549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd153550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd153551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd153552: begin  
rid<=0;
end
18'd153601: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=14;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16506;
 end   
18'd153602: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=78;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd153603: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=68;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd153604: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=33;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd153605: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=20;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd153606: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=91;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd153607: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd153608: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd153609: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd153610: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd153611: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd153612: begin  
  clrr<=0;
  maplen<=6;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd153742: begin  
rid<=1;
end
18'd153743: begin  
end
18'd153744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd153745: begin  
rid<=0;
end
18'd153801: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=89;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6942;
 end   
18'd153802: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=98;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7654;
 end   
18'd153803: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=16;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1268;
 end   
18'd153804: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=30;
 end   
18'd153805: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=57;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=4486;
 end   
18'd153806: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=32;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=2546;
 end   
18'd153807: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=3;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=294;
 end   
18'd153808: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=62;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=4906;
 end   
18'd153809: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=82;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=6476;
 end   
18'd153810: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd153942: begin  
rid<=1;
end
18'd153943: begin  
end
18'd153944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd153945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd153946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd153947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd153948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd153949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd153950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd153951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd153952: begin  
check<=expctdoutput[8]-outcheck;
end
18'd153953: begin  
rid<=0;
end
18'd154001: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=74;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=21104;
 end   
18'd154002: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=69;
   mapp<=61;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=21932;
 end   
18'd154003: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=99;
   mapp<=25;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=17159;
 end   
18'd154004: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=97;
   mapp<=84;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=19683;
 end   
18'd154005: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=98;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd154006: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=34;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd154007: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd154008: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd154009: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd154010: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd154011: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd154012: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd154013: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21104;
 end   
18'd154014: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21104;
 end   
18'd154015: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21104;
 end   
18'd154142: begin  
rid<=1;
end
18'd154143: begin  
end
18'd154144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd154145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd154146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd154147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd154148: begin  
rid<=0;
end
18'd154201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=80;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=21895;
 end   
18'd154202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=91;
   mapp<=88;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=18641;
 end   
18'd154203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=61;
   mapp<=51;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=17565;
 end   
18'd154204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=88;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd154205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=39;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd154206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=60;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd154207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd154208: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd154209: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd154210: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd154342: begin  
rid<=1;
end
18'd154343: begin  
end
18'd154344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd154345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd154346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd154347: begin  
rid<=0;
end
18'd154401: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=21;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=231;
 end   
18'd154402: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=33;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=703;
 end   
18'd154403: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=26;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=566;
 end   
18'd154404: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=52;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=1122;
 end   
18'd154405: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=46;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=1006;
 end   
18'd154406: begin  
  clrr<=0;
  maplen<=5;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd154542: begin  
rid<=1;
end
18'd154543: begin  
end
18'd154544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd154545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd154546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd154547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd154548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd154549: begin  
rid<=0;
end
18'd154601: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=67;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=20025;
 end   
18'd154602: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=98;
   mapp<=45;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=18326;
 end   
18'd154603: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=57;
   mapp<=25;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=17622;
 end   
18'd154604: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=41;
   mapp<=23;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=20679;
 end   
18'd154605: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=50;
   mapp<=76;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=21349;
 end   
18'd154606: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=52;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd154607: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=49;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd154608: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd154609: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd154610: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd154611: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd154612: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd154613: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20025;
 end   
18'd154614: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20025;
 end   
18'd154615: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20025;
 end   
18'd154616: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20025;
 end   
18'd154617: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20025;
 end   
18'd154618: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20025;
 end   
18'd154742: begin  
rid<=1;
end
18'd154743: begin  
end
18'd154744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd154745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd154746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd154747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd154748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd154749: begin  
rid<=0;
end
18'd154801: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=13;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6810;
 end   
18'd154802: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=49;
   mapp<=14;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10691;
 end   
18'd154803: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=24;
   mapp<=53;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=7633;
 end   
18'd154804: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=42;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd154805: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=54;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd154806: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=17;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd154807: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=40;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd154808: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd154809: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd154810: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd154811: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd154812: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd154813: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6810;
 end   
18'd154814: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6810;
 end   
18'd154815: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6810;
 end   
18'd154816: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6810;
 end   
18'd154942: begin  
rid<=1;
end
18'd154943: begin  
end
18'd154944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd154945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd154946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd154947: begin  
rid<=0;
end
18'd155001: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=97;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12607;
 end   
18'd155002: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=87;
   mapp<=28;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=12400;
 end   
18'd155003: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=0;
   mapp<=63;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=7531;
 end   
18'd155004: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=86;
   mapp<=63;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=8976;
 end   
18'd155005: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=43;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=5605;
 end   
18'd155006: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=38;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=4432;
 end   
18'd155007: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=18;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=8369;
 end   
18'd155008: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=20;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd155009: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd155010: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=97;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd155011: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd155012: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd155013: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12607;
 end   
18'd155014: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12607;
 end   
18'd155142: begin  
rid<=1;
end
18'd155143: begin  
end
18'd155144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd155145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd155146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd155147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd155148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd155149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd155150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd155151: begin  
rid<=0;
end
18'd155201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=35;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13004;
 end   
18'd155202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=90;
   mapp<=70;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=18214;
 end   
18'd155203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=97;
   mapp<=37;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=15722;
 end   
18'd155204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=92;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=9519;
 end   
18'd155205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=17;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd155206: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=3;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd155207: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd155208: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd155209: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd155342: begin  
rid<=1;
end
18'd155343: begin  
end
18'd155344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd155345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd155346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd155347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd155348: begin  
rid<=0;
end
18'd155401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=98;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=20712;
 end   
18'd155402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=50;
   mapp<=19;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=19062;
 end   
18'd155403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=90;
   mapp<=97;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=24410;
 end   
18'd155404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=48;
   mapp<=54;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=21094;
 end   
18'd155405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=56;
   mapp<=28;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=18906;
 end   
18'd155406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=24;
   mapp<=74;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=21166;
 end   
18'd155407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd155408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd155409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd155410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd155411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd155412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd155413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20712;
 end   
18'd155414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20712;
 end   
18'd155415: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20712;
 end   
18'd155416: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20712;
 end   
18'd155417: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=20712;
 end   
18'd155542: begin  
rid<=1;
end
18'd155543: begin  
end
18'd155544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd155545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd155546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd155547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd155548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd155549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd155550: begin  
rid<=0;
end
18'd155601: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=85;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=425;
 end   
18'd155602: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5790;
 end   
18'd155603: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=40;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=3420;
 end   
18'd155604: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=87;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=7425;
 end   
18'd155605: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=55;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=4715;
 end   
18'd155606: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=28;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=2430;
 end   
18'd155607: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=55;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=4735;
 end   
18'd155608: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd155609: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd155610: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd155742: begin  
rid<=1;
end
18'd155743: begin  
end
18'd155744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd155745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd155746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd155747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd155748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd155749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd155750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd155751: begin  
rid<=0;
end
18'd155801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=10;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11397;
 end   
18'd155802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=47;
   mapp<=75;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=16241;
 end   
18'd155803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=81;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd155804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=55;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd155805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=74;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd155806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=38;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd155807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd155808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd155809: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd155810: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd155811: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd155812: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd155813: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11397;
 end   
18'd155942: begin  
rid<=1;
end
18'd155943: begin  
end
18'd155944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd155945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd155946: begin  
rid<=0;
end
18'd156001: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=74;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9604;
 end   
18'd156002: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=69;
   mapp<=15;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=14229;
 end   
18'd156003: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=52;
   mapp<=12;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=13138;
 end   
18'd156004: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=16;
   mapp<=97;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=16194;
 end   
18'd156005: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=64;
   mapp<=31;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=14081;
 end   
18'd156006: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=59;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd156007: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=86;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd156008: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=51;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd156009: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=87;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd156010: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=72;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd156011: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=45;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd156012: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd156013: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9604;
 end   
18'd156014: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9604;
 end   
18'd156015: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9604;
 end   
18'd156016: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9604;
 end   
18'd156017: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9604;
 end   
18'd156018: begin  
  clrr<=0;
  maplen<=7;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9604;
 end   
18'd156142: begin  
rid<=1;
end
18'd156143: begin  
end
18'd156144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd156145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd156146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd156147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd156148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd156149: begin  
rid<=0;
end
18'd156201: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=57;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=291;
 end   
18'd156202: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=18;
   mapp<=13;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2353;
 end   
18'd156203: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=89;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=5669;
 end   
18'd156204: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=32;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=3438;
 end   
18'd156205: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=88;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=5272;
 end   
18'd156206: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=12;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=1436;
 end   
18'd156207: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=39;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=3903;
 end   
18'd156208: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd156209: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd156210: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd156342: begin  
rid<=1;
end
18'd156343: begin  
end
18'd156344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd156345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd156346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd156347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd156348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd156349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd156350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd156351: begin  
rid<=0;
end
18'd156401: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=71;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=17019;
 end   
18'd156402: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=6;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=20278;
 end   
18'd156403: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=52;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd156404: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=86;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd156405: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=44;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd156406: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=40;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd156407: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd156408: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd156409: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd156410: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd156411: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd156412: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd156413: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17019;
 end   
18'd156542: begin  
rid<=1;
end
18'd156543: begin  
end
18'd156544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd156545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd156546: begin  
rid<=0;
end
18'd156601: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=98;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15516;
 end   
18'd156602: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=87;
   mapp<=73;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10374;
 end   
18'd156603: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=21;
   mapp<=59;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=4477;
 end   
18'd156604: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=2;
   mapp<=92;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=6916;
 end   
18'd156605: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=20;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=7585;
 end   
18'd156606: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=16;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=8343;
 end   
18'd156607: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=47;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=7038;
 end   
18'd156608: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=22;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=5591;
 end   
18'd156609: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=25;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd156610: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=2;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd156611: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=20;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd156612: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd156613: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15516;
 end   
18'd156614: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15516;
 end   
18'd156615: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15516;
 end   
18'd156742: begin  
rid<=1;
end
18'd156743: begin  
end
18'd156744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd156745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd156746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd156747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd156748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd156749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd156750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd156751: begin  
check<=expctdoutput[7]-outcheck;
end
18'd156752: begin  
rid<=0;
end
18'd156801: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=68;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9036;
 end   
18'd156802: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=38;
   mapp<=69;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9916;
 end   
18'd156803: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=74;
   mapp<=83;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5591;
 end   
18'd156804: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=56;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd156805: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=17;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd156806: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd156807: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd156808: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd156942: begin  
rid<=1;
end
18'd156943: begin  
end
18'd156944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd156945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd156946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd156947: begin  
rid<=0;
end
18'd157001: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=48;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1536;
 end   
18'd157002: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=47;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1514;
 end   
18'd157003: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=44;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1428;
 end   
18'd157004: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=9;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=318;
 end   
18'd157005: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=46;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=1512;
 end   
18'd157006: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=56;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=1842;
 end   
18'd157007: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=70;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=2300;
 end   
18'd157008: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=41;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=1382;
 end   
18'd157009: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=39;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=1328;
 end   
18'd157010: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd157142: begin  
rid<=1;
end
18'd157143: begin  
end
18'd157144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd157145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd157146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd157147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd157148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd157149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd157150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd157151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd157152: begin  
check<=expctdoutput[8]-outcheck;
end
18'd157153: begin  
rid<=0;
end
18'd157201: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=28;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3911;
 end   
18'd157202: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=88;
   mapp<=31;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5534;
 end   
18'd157203: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=39;
   mapp<=21;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=10688;
 end   
18'd157204: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd157205: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd157206: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd157207: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd157208: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd157342: begin  
rid<=1;
end
18'd157343: begin  
end
18'd157344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd157345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd157346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd157347: begin  
rid<=0;
end
18'd157401: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=84;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4620;
 end   
18'd157402: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=58;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3200;
 end   
18'd157403: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=84;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=4640;
 end   
18'd157404: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd157542: begin  
rid<=1;
end
18'd157543: begin  
end
18'd157544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd157545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd157546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd157547: begin  
rid<=0;
end
18'd157601: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=71;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6319;
 end   
18'd157602: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=94;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8376;
 end   
18'd157603: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=85;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=7585;
 end   
18'd157604: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd157742: begin  
rid<=1;
end
18'd157743: begin  
end
18'd157744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd157745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd157746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd157747: begin  
rid<=0;
end
18'd157801: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=54;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4050;
 end   
18'd157802: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=61;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=3304;
 end   
18'd157803: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=24;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=1316;
 end   
18'd157804: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=71;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=3864;
 end   
18'd157805: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=66;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=3604;
 end   
18'd157806: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=35;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=1940;
 end   
18'd157807: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=59;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=3246;
 end   
18'd157808: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=40;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=2230;
 end   
18'd157809: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=43;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=2402;
 end   
18'd157810: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=56;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[9]<=3114;
 end   
18'd157811: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd157942: begin  
rid<=1;
end
18'd157943: begin  
end
18'd157944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd157945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd157946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd157947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd157948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd157949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd157950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd157951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd157952: begin  
check<=expctdoutput[8]-outcheck;
end
18'd157953: begin  
check<=expctdoutput[9]-outcheck;
end
18'd157954: begin  
rid<=0;
end
18'd158001: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=23;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2392;
 end   
18'd158002: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=37;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd158003: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=38;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd158004: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd158005: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd158006: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd158142: begin  
rid<=1;
end
18'd158143: begin  
end
18'd158144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd158145: begin  
rid<=0;
end
18'd158201: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=2;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=182;
 end   
18'd158202: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=89;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8109;
 end   
18'd158203: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=87;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=7937;
 end   
18'd158204: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=97;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=8857;
 end   
18'd158205: begin  
  clrr<=0;
  maplen<=1;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd158342: begin  
rid<=1;
end
18'd158343: begin  
end
18'd158344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd158345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd158346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd158347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd158348: begin  
rid<=0;
end
18'd158401: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=12;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=18343;
 end   
18'd158402: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=98;
   mapp<=26;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=17404;
 end   
18'd158403: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=72;
   mapp<=23;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=24526;
 end   
18'd158404: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=55;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd158405: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=71;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd158406: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=9;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd158407: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=53;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd158408: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd158409: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd158410: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd158411: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd158412: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd158413: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18343;
 end   
18'd158414: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18343;
 end   
18'd158415: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18343;
 end   
18'd158416: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18343;
 end   
18'd158542: begin  
rid<=1;
end
18'd158543: begin  
end
18'd158544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd158545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd158546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd158547: begin  
rid<=0;
end
18'd158601: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=4;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1667;
 end   
18'd158602: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=18;
   mapp<=12;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4095;
 end   
18'd158603: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=45;
   mapp<=16;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6290;
 end   
18'd158604: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=13;
   mapp<=55;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=5545;
 end   
18'd158605: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=98;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=5361;
 end   
18'd158606: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=62;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=5878;
 end   
18'd158607: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=57;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=3658;
 end   
18'd158608: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd158609: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd158610: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd158611: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd158612: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd158613: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=1667;
 end   
18'd158614: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=1667;
 end   
18'd158742: begin  
rid<=1;
end
18'd158743: begin  
end
18'd158744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd158745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd158746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd158747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd158748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd158749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd158750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd158751: begin  
rid<=0;
end
18'd158801: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=60;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1980;
 end   
18'd158802: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=54;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=3250;
 end   
18'd158803: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=18;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=1100;
 end   
18'd158804: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=30;
 end   
18'd158805: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=29;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=1780;
 end   
18'd158806: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=61;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=3710;
 end   
18'd158807: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=32;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=1980;
 end   
18'd158808: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=58;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=3550;
 end   
18'd158809: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=46;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=2840;
 end   
18'd158810: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd158942: begin  
rid<=1;
end
18'd158943: begin  
end
18'd158944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd158945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd158946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd158947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd158948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd158949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd158950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd158951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd158952: begin  
check<=expctdoutput[8]-outcheck;
end
18'd158953: begin  
rid<=0;
end
18'd159001: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=31;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1049;
 end   
18'd159002: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=39;
   mapp<=12;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=961;
 end   
18'd159003: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=9;
   mapp<=6;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1073;
 end   
18'd159004: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=30;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=1842;
 end   
18'd159005: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=90;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd159006: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd159007: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd159008: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd159009: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd159142: begin  
rid<=1;
end
18'd159143: begin  
end
18'd159144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd159145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd159146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd159147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd159148: begin  
rid<=0;
end
18'd159201: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=78;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=25153;
 end   
18'd159202: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=56;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd159203: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=34;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd159204: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=74;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd159205: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=47;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd159206: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=95;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd159207: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd159208: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=61;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd159209: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=63;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd159210: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd159211: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd159212: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd159213: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25153;
 end   
18'd159214: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25153;
 end   
18'd159215: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25153;
 end   
18'd159216: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25153;
 end   
18'd159217: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25153;
 end   
18'd159218: begin  
  clrr<=0;
  maplen<=9;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25153;
 end   
18'd159342: begin  
rid<=1;
end
18'd159343: begin  
end
18'd159344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd159345: begin  
rid<=0;
end
18'd159401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=12;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=23429;
 end   
18'd159402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=92;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=17669;
 end   
18'd159403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=84;
   mapp<=26;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=22765;
 end   
18'd159404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=36;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd159405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=61;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd159406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=2;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd159407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=99;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd159408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=17;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd159409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=9;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd159410: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=52;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd159411: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd159412: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd159413: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23429;
 end   
18'd159414: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23429;
 end   
18'd159415: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23429;
 end   
18'd159416: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23429;
 end   
18'd159417: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23429;
 end   
18'd159418: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23429;
 end   
18'd159542: begin  
rid<=1;
end
18'd159543: begin  
end
18'd159544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd159545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd159546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd159547: begin  
rid<=0;
end
18'd159601: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=63;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9760;
 end   
18'd159602: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=73;
   mapp<=66;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9371;
 end   
18'd159603: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=31;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6354;
 end   
18'd159604: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=3;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=5381;
 end   
18'd159605: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=55;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=6888;
 end   
18'd159606: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=37;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=6684;
 end   
18'd159607: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=22;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=10184;
 end   
18'd159608: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=87;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=11451;
 end   
18'd159609: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd159610: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd159611: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd159612: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd159613: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9760;
 end   
18'd159742: begin  
rid<=1;
end
18'd159743: begin  
end
18'd159744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd159745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd159746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd159747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd159748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd159749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd159750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd159751: begin  
check<=expctdoutput[7]-outcheck;
end
18'd159752: begin  
rid<=0;
end
18'd159801: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=35;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16760;
 end   
18'd159802: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=97;
   mapp<=58;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=19945;
 end   
18'd159803: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=25;
   mapp<=92;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12742;
 end   
18'd159804: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=7;
   mapp<=63;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=14461;
 end   
18'd159805: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=84;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd159806: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd159807: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd159808: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd159809: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd159810: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd159811: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd159812: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd159813: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16760;
 end   
18'd159942: begin  
rid<=1;
end
18'd159943: begin  
end
18'd159944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd159945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd159946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd159947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd159948: begin  
rid<=0;
end
18'd160001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=29;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16186;
 end   
18'd160002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=93;
   mapp<=94;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=19263;
 end   
18'd160003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=47;
   mapp<=73;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12350;
 end   
18'd160004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=61;
   mapp<=4;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=12426;
 end   
18'd160005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=28;
   mapp<=59;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=9674;
 end   
18'd160006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=59;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=10889;
 end   
18'd160007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=15;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=7676;
 end   
18'd160008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd160009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=15;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd160010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=66;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd160011: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd160012: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd160013: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16186;
 end   
18'd160014: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16186;
 end   
18'd160015: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16186;
 end   
18'd160016: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16186;
 end   
18'd160142: begin  
rid<=1;
end
18'd160143: begin  
end
18'd160144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd160145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd160146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd160147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd160148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd160149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd160150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd160151: begin  
rid<=0;
end
18'd160201: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=79;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10470;
 end   
18'd160202: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=88;
   mapp<=31;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10897;
 end   
18'd160203: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=73;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8600;
 end   
18'd160204: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=46;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=7297;
 end   
18'd160205: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=89;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=11242;
 end   
18'd160206: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=80;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=10401;
 end   
18'd160207: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=81;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=7998;
 end   
18'd160208: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=2550;
 end   
18'd160209: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=80;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=10617;
 end   
18'd160210: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=87;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[9]<=9887;
 end   
18'd160211: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=41;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd160212: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd160213: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10470;
 end   
18'd160342: begin  
rid<=1;
end
18'd160343: begin  
end
18'd160344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd160345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd160346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd160347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd160348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd160349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd160350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd160351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd160352: begin  
check<=expctdoutput[8]-outcheck;
end
18'd160353: begin  
check<=expctdoutput[9]-outcheck;
end
18'd160354: begin  
rid<=0;
end
18'd160401: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=73;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7866;
 end   
18'd160402: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=8;
   mapp<=89;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1595;
 end   
18'd160403: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=9;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5352;
 end   
18'd160404: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=50;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=5642;
 end   
18'd160405: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=8;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd160406: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd160407: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd160542: begin  
rid<=1;
end
18'd160543: begin  
end
18'd160544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd160545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd160546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd160547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd160548: begin  
rid<=0;
end
18'd160601: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=50;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1250;
 end   
18'd160602: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=4;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=110;
 end   
18'd160603: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=36;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=920;
 end   
18'd160604: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=67;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=1705;
 end   
18'd160605: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=54;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=1390;
 end   
18'd160606: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=85;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=2175;
 end   
18'd160607: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=85;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=2185;
 end   
18'd160608: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=21;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=595;
 end   
18'd160609: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=28;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=780;
 end   
18'd160610: begin  
  clrr<=0;
  maplen<=1;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd160742: begin  
rid<=1;
end
18'd160743: begin  
end
18'd160744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd160745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd160746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd160747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd160748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd160749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd160750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd160751: begin  
check<=expctdoutput[7]-outcheck;
end
18'd160752: begin  
check<=expctdoutput[8]-outcheck;
end
18'd160753: begin  
rid<=0;
end
18'd160801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=48;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15547;
 end   
18'd160802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=56;
   mapp<=44;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=18377;
 end   
18'd160803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=31;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd160804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=41;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd160805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=78;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd160806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=73;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd160807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=89;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd160808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=97;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd160809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd160810: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd160811: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd160812: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd160813: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15547;
 end   
18'd160814: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15547;
 end   
18'd160815: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15547;
 end   
18'd160942: begin  
rid<=1;
end
18'd160943: begin  
end
18'd160944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd160945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd160946: begin  
rid<=0;
end
18'd161001: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=89;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9036;
 end   
18'd161002: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=98;
   mapp<=25;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8605;
 end   
18'd161003: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=65;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=8647;
 end   
18'd161004: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=29;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=7511;
 end   
18'd161005: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=50;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=8018;
 end   
18'd161006: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd161007: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd161008: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd161142: begin  
rid<=1;
end
18'd161143: begin  
end
18'd161144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd161145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd161146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd161147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd161148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd161149: begin  
rid<=0;
end
18'd161201: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=22;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9386;
 end   
18'd161202: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=16;
   mapp<=39;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5493;
 end   
18'd161203: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=22;
   mapp<=37;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5339;
 end   
18'd161204: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=25;
   mapp<=34;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=9875;
 end   
18'd161205: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=79;
   mapp<=84;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=12134;
 end   
18'd161206: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=15;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=8289;
 end   
18'd161207: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd161208: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd161209: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd161210: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd161211: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd161212: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd161213: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9386;
 end   
18'd161214: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9386;
 end   
18'd161215: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9386;
 end   
18'd161342: begin  
rid<=1;
end
18'd161343: begin  
end
18'd161344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd161345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd161346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd161347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd161348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd161349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd161350: begin  
rid<=0;
end
18'd161401: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=18;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1637;
 end   
18'd161402: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=20;
   mapp<=4;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6592;
 end   
18'd161403: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=3;
   mapp<=93;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8105;
 end   
18'd161404: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=75;
   mapp<=0;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=8269;
 end   
18'd161405: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=62;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=9761;
 end   
18'd161406: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=83;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=4886;
 end   
18'd161407: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=90;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=10336;
 end   
18'd161408: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd161409: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd161410: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd161411: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd161412: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd161413: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=1637;
 end   
18'd161414: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=1637;
 end   
18'd161542: begin  
rid<=1;
end
18'd161543: begin  
end
18'd161544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd161545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd161546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd161547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd161548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd161549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd161550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd161551: begin  
rid<=0;
end
18'd161601: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=87;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9358;
 end   
18'd161602: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=16;
   mapp<=8;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5054;
 end   
18'd161603: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=18;
   mapp<=41;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12757;
 end   
18'd161604: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=18;
   mapp<=98;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=11460;
 end   
18'd161605: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=68;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd161606: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd161607: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd161608: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd161609: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd161610: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd161611: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd161612: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd161613: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9358;
 end   
18'd161742: begin  
rid<=1;
end
18'd161743: begin  
end
18'd161744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd161745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd161746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd161747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd161748: begin  
rid<=0;
end
18'd161801: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=10;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4498;
 end   
18'd161802: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=44;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4192;
 end   
18'd161803: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=73;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=3038;
 end   
18'd161804: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=52;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=1210;
 end   
18'd161805: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=15;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=2654;
 end   
18'd161806: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=56;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=1842;
 end   
18'd161807: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=28;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=1000;
 end   
18'd161808: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=15;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=1056;
 end   
18'd161809: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=19;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=2162;
 end   
18'd161810: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=43;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[9]<=2632;
 end   
18'd161811: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd161812: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd161813: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=4498;
 end   
18'd161942: begin  
rid<=1;
end
18'd161943: begin  
end
18'd161944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd161945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd161946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd161947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd161948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd161949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd161950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd161951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd161952: begin  
check<=expctdoutput[8]-outcheck;
end
18'd161953: begin  
check<=expctdoutput[9]-outcheck;
end
18'd161954: begin  
rid<=0;
end
18'd162001: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=35;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6480;
 end   
18'd162002: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=4;
   mapp<=37;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4692;
 end   
18'd162003: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=32;
   mapp<=12;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8444;
 end   
18'd162004: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=16;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd162005: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=91;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd162006: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd162007: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd162008: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd162009: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd162010: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd162011: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd162012: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd162142: begin  
rid<=1;
end
18'd162143: begin  
end
18'd162144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd162145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd162146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd162147: begin  
rid<=0;
end
18'd162201: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=89;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5292;
 end   
18'd162202: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=25;
   mapp<=23;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4007;
 end   
18'd162203: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=78;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=7787;
 end   
18'd162204: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=33;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=4517;
 end   
18'd162205: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=62;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=7808;
 end   
18'd162206: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=90;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=8760;
 end   
18'd162207: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=28;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=3152;
 end   
18'd162208: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=24;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=4231;
 end   
18'd162209: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd162210: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd162211: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd162342: begin  
rid<=1;
end
18'd162343: begin  
end
18'd162344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd162345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd162346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd162347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd162348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd162349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd162350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd162351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd162352: begin  
rid<=0;
end
18'd162401: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=67;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15922;
 end   
18'd162402: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=37;
   mapp<=96;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=17087;
 end   
18'd162403: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=55;
   mapp<=62;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=19108;
 end   
18'd162404: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=75;
   mapp<=63;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=18248;
 end   
18'd162405: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=54;
   mapp<=35;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=18541;
 end   
18'd162406: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=70;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=16797;
 end   
18'd162407: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=63;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=16229;
 end   
18'd162408: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=60;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd162409: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=63;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd162410: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd162411: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=94;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd162412: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd162413: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15922;
 end   
18'd162414: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15922;
 end   
18'd162415: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15922;
 end   
18'd162416: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15922;
 end   
18'd162542: begin  
rid<=1;
end
18'd162543: begin  
end
18'd162544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd162545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd162546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd162547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd162548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd162549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd162550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd162551: begin  
rid<=0;
end
18'd162601: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=64;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=576;
 end   
18'd162602: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=12;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=118;
 end   
18'd162603: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=24;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=236;
 end   
18'd162604: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=34;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=336;
 end   
18'd162605: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=6;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=94;
 end   
18'd162606: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=81;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=779;
 end   
18'd162607: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=90;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=870;
 end   
18'd162608: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=34;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=376;
 end   
18'd162609: begin  
  clrr<=0;
  maplen<=1;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd162742: begin  
rid<=1;
end
18'd162743: begin  
end
18'd162744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd162745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd162746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd162747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd162748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd162749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd162750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd162751: begin  
check<=expctdoutput[7]-outcheck;
end
18'd162752: begin  
rid<=0;
end
18'd162801: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=50;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6424;
 end   
18'd162802: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=44;
   mapp<=19;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8558;
 end   
18'd162803: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=18;
   mapp<=26;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=4890;
 end   
18'd162804: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=16;
   mapp<=70;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=3461;
 end   
18'd162805: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=61;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=7314;
 end   
18'd162806: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=22;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=2810;
 end   
18'd162807: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=6;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=3842;
 end   
18'd162808: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=26;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd162809: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=3;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd162810: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=39;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd162811: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd162812: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd162813: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6424;
 end   
18'd162814: begin  
  clrr<=0;
  maplen<=4;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6424;
 end   
18'd162942: begin  
rid<=1;
end
18'd162943: begin  
end
18'd162944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd162945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd162946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd162947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd162948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd162949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd162950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd162951: begin  
rid<=0;
end
18'd163001: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=32;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1632;
 end   
18'd163002: begin  
  clrr<=0;
  maplen<=1;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd163142: begin  
rid<=1;
end
18'd163143: begin  
end
18'd163144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd163145: begin  
rid<=0;
end
18'd163201: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=34;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7566;
 end   
18'd163202: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=51;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7624;
 end   
18'd163203: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=40;
   mapp<=2;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=13369;
 end   
18'd163204: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=10;
   mapp<=63;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=14946;
 end   
18'd163205: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=38;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd163206: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=7;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd163207: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=49;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd163208: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=51;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd163209: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd163210: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd163211: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd163212: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd163213: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7566;
 end   
18'd163214: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7566;
 end   
18'd163215: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7566;
 end   
18'd163216: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7566;
 end   
18'd163217: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7566;
 end   
18'd163218: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7566;
 end   
18'd163219: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7566;
 end   
18'd163342: begin  
rid<=1;
end
18'd163343: begin  
end
18'd163344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd163345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd163346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd163347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd163348: begin  
rid<=0;
end
18'd163401: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=73;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=29293;
 end   
18'd163402: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=89;
   mapp<=71;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=25623;
 end   
18'd163403: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=85;
   mapp<=21;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=27232;
 end   
18'd163404: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=81;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd163405: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=55;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd163406: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=87;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd163407: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=94;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd163408: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=6;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd163409: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd163410: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd163411: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd163412: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd163413: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29293;
 end   
18'd163414: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29293;
 end   
18'd163415: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29293;
 end   
18'd163416: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29293;
 end   
18'd163417: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29293;
 end   
18'd163418: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29293;
 end   
18'd163542: begin  
rid<=1;
end
18'd163543: begin  
end
18'd163544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd163545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd163546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd163547: begin  
rid<=0;
end
18'd163601: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=71;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13857;
 end   
18'd163602: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=52;
   mapp<=87;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11891;
 end   
18'd163603: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=95;
   mapp<=42;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=13868;
 end   
18'd163604: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=21;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd163605: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=1;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd163606: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=87;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd163607: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd163608: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd163609: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd163610: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd163742: begin  
rid<=1;
end
18'd163743: begin  
end
18'd163744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd163745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd163746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd163747: begin  
rid<=0;
end
18'd163801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=72;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4791;
 end   
18'd163802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=21;
   mapp<=91;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7192;
 end   
18'd163803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=30;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=3377;
 end   
18'd163804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=57;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=5205;
 end   
18'd163805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=51;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=3796;
 end   
18'd163806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd163807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd163808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd163942: begin  
rid<=1;
end
18'd163943: begin  
end
18'd163944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd163945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd163946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd163947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd163948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd163949: begin  
rid<=0;
end
18'd164001: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=22;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4484;
 end   
18'd164002: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=78;
   mapp<=51;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7216;
 end   
18'd164003: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=78;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=9380;
 end   
18'd164004: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=98;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=8894;
 end   
18'd164005: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=86;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=8796;
 end   
18'd164006: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=88;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=3624;
 end   
18'd164007: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=21;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=1380;
 end   
18'd164008: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=11;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=312;
 end   
18'd164009: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=2264;
 end   
18'd164010: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=28;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[9]<=1408;
 end   
18'd164011: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=9;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd164012: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd164013: begin  
  clrr<=0;
  maplen<=11;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=4484;
 end   
18'd164142: begin  
rid<=1;
end
18'd164143: begin  
end
18'd164144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd164145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd164146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd164147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd164148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd164149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd164150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd164151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd164152: begin  
check<=expctdoutput[8]-outcheck;
end
18'd164153: begin  
check<=expctdoutput[9]-outcheck;
end
18'd164154: begin  
rid<=0;
end
18'd164201: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=50;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16336;
 end   
18'd164202: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=86;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=15231;
 end   
18'd164203: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=7;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd164204: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=26;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd164205: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=49;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd164206: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=73;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd164207: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=64;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd164208: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd164209: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd164210: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd164211: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd164212: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd164213: begin  
  clrr<=0;
  maplen<=6;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16336;
 end   
18'd164342: begin  
rid<=1;
end
18'd164343: begin  
end
18'd164344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd164345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd164346: begin  
rid<=0;
end
18'd164401: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=70;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12250;
 end   
18'd164402: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=53;
   mapp<=22;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9688;
 end   
18'd164403: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=4;
   mapp<=46;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=10262;
 end   
18'd164404: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=56;
   mapp<=46;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=9405;
 end   
18'd164405: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=54;
   mapp<=31;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=10200;
 end   
18'd164406: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=70;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=9386;
 end   
18'd164407: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd164408: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd164409: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd164410: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd164411: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd164412: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd164413: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12250;
 end   
18'd164414: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12250;
 end   
18'd164415: begin  
  clrr<=0;
  maplen<=10;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12250;
 end   
18'd164542: begin  
rid<=1;
end
18'd164543: begin  
end
18'd164544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd164545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd164546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd164547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd164548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd164549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd164550: begin  
rid<=0;
end
18'd164601: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=93;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9596;
 end   
18'd164602: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=91;
   mapp<=19;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8227;
 end   
18'd164603: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=40;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd164604: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=57;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd164605: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=0;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd164606: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd164607: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd164608: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd164609: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd164742: begin  
rid<=1;
end
18'd164743: begin  
end
18'd164744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd164745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd164746: begin  
rid<=0;
end
18'd164801: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=7;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11164;
 end   
18'd164802: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=51;
   mapp<=31;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11113;
 end   
18'd164803: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=22;
   mapp<=6;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12663;
 end   
18'd164804: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=4;
   mapp<=88;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=8185;
 end   
18'd164805: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=90;
   mapp<=55;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=12667;
 end   
18'd164806: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=81;
   mapp<=45;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=19303;
 end   
18'd164807: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd164808: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd164809: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd164810: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd164811: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd164812: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd164813: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11164;
 end   
18'd164814: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11164;
 end   
18'd164815: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11164;
 end   
18'd164816: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11164;
 end   
18'd164817: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11164;
 end   
18'd164942: begin  
rid<=1;
end
18'd164943: begin  
end
18'd164944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd164945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd164946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd164947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd164948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd164949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd164950: begin  
rid<=0;
end
18'd165001: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=14;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3054;
 end   
18'd165002: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=64;
   mapp<=44;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1394;
 end   
18'd165003: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd165004: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd165005: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd165142: begin  
rid<=1;
end
18'd165143: begin  
end
18'd165144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd165145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd165146: begin  
rid<=0;
end
18'd165201: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=86;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9577;
 end   
18'd165202: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=79;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd165203: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd165204: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd165342: begin  
rid<=1;
end
18'd165343: begin  
end
18'd165344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd165345: begin  
rid<=0;
end
18'd165401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=84;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=21814;
 end   
18'd165402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=58;
   mapp<=82;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=24445;
 end   
18'd165403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=4;
   mapp<=39;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=19006;
 end   
18'd165404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=48;
   mapp<=27;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=15853;
 end   
18'd165405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=58;
   mapp<=66;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=18319;
 end   
18'd165406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=83;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd165407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=52;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd165408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd165409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd165410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd165411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd165412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd165413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21814;
 end   
18'd165414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21814;
 end   
18'd165415: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21814;
 end   
18'd165416: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21814;
 end   
18'd165417: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21814;
 end   
18'd165418: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21814;
 end   
18'd165542: begin  
rid<=1;
end
18'd165543: begin  
end
18'd165544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd165545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd165546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd165547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd165548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd165549: begin  
rid<=0;
end
18'd165601: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=55;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13427;
 end   
18'd165602: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=39;
   mapp<=74;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=15827;
 end   
18'd165603: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=53;
   mapp<=22;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12113;
 end   
18'd165604: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=76;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd165605: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd165606: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd165607: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd165608: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd165609: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd165610: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd165742: begin  
rid<=1;
end
18'd165743: begin  
end
18'd165744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd165745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd165746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd165747: begin  
rid<=0;
end
18'd165801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=10;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14238;
 end   
18'd165802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=80;
   mapp<=82;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13015;
 end   
18'd165803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=60;
   mapp<=31;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=14228;
 end   
18'd165804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=78;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd165805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=27;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd165806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd165807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd165808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd165809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd165810: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd165811: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd165812: begin  
  clrr<=0;
  maplen<=7;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd165942: begin  
rid<=1;
end
18'd165943: begin  
end
18'd165944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd165945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd165946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd165947: begin  
rid<=0;
end
18'd166001: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=15;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8380;
 end   
18'd166002: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=71;
   mapp<=30;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=18592;
 end   
18'd166003: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=29;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd166004: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=6;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd166005: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=1;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd166006: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=94;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd166007: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=84;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd166008: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=15;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd166009: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=67;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd166010: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd166011: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd166012: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd166013: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8380;
 end   
18'd166014: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8380;
 end   
18'd166015: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8380;
 end   
18'd166016: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8380;
 end   
18'd166017: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8380;
 end   
18'd166142: begin  
rid<=1;
end
18'd166143: begin  
end
18'd166144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd166145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd166146: begin  
rid<=0;
end
18'd166201: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=82;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7842;
 end   
18'd166202: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=26;
   mapp<=84;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6676;
 end   
18'd166203: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=58;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=4946;
 end   
18'd166204: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=11;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=1125;
 end   
18'd166205: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=4;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=4096;
 end   
18'd166206: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=45;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=7523;
 end   
18'd166207: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=52;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=10452;
 end   
18'd166208: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=81;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=8431;
 end   
18'd166209: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=33;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd166210: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd166211: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd166342: begin  
rid<=1;
end
18'd166343: begin  
end
18'd166344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd166345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd166346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd166347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd166348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd166349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd166350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd166351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd166352: begin  
rid<=0;
end
18'd166401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=33;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=17246;
 end   
18'd166402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=54;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd166403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=49;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd166404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=6;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd166405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=4;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd166406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=29;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd166407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=95;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd166408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=66;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd166409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd166410: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd166411: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd166412: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd166413: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17246;
 end   
18'd166414: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17246;
 end   
18'd166415: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17246;
 end   
18'd166416: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17246;
 end   
18'd166542: begin  
rid<=1;
end
18'd166543: begin  
end
18'd166544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd166545: begin  
rid<=0;
end
18'd166601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=62;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1686;
 end   
18'd166602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=34;
   mapp<=4;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1754;
 end   
18'd166603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=44;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=2952;
 end   
18'd166604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=6;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=3768;
 end   
18'd166605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=99;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=7606;
 end   
18'd166606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=42;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=5986;
 end   
18'd166607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=98;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=7870;
 end   
18'd166608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=51;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=4388;
 end   
18'd166609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd166610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd166611: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd166742: begin  
rid<=1;
end
18'd166743: begin  
end
18'd166744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd166745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd166746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd166747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd166748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd166749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd166750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd166751: begin  
check<=expctdoutput[7]-outcheck;
end
18'd166752: begin  
rid<=0;
end
18'd166801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=73;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16140;
 end   
18'd166802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=79;
   mapp<=97;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=14830;
 end   
18'd166803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=55;
   mapp<=36;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12099;
 end   
18'd166804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=89;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=12808;
 end   
18'd166805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=44;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=10801;
 end   
18'd166806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd166807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd166808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd166809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd166810: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd166942: begin  
rid<=1;
end
18'd166943: begin  
end
18'd166944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd166945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd166946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd166947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd166948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd166949: begin  
rid<=0;
end
18'd167001: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=35;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=23623;
 end   
18'd167002: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=71;
   mapp<=25;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=19969;
 end   
18'd167003: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=63;
   mapp<=50;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=22634;
 end   
18'd167004: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=54;
   mapp<=86;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=18790;
 end   
18'd167005: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=88;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd167006: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=30;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd167007: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=66;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd167008: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd167009: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd167010: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd167011: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd167012: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd167013: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23623;
 end   
18'd167014: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23623;
 end   
18'd167015: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23623;
 end   
18'd167016: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23623;
 end   
18'd167017: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23623;
 end   
18'd167142: begin  
rid<=1;
end
18'd167143: begin  
end
18'd167144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd167145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd167146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd167147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd167148: begin  
rid<=0;
end
18'd167201: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=34;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8878;
 end   
18'd167202: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=96;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11884;
 end   
18'd167203: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=67;
   mapp<=84;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12584;
 end   
18'd167204: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=2;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd167205: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd167206: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd167207: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd167208: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd167209: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd167210: begin  
  clrr<=0;
  maplen<=6;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd167342: begin  
rid<=1;
end
18'd167343: begin  
end
18'd167344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd167345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd167346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd167347: begin  
rid<=0;
end
18'd167401: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=35;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7900;
 end   
18'd167402: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=78;
   mapp<=88;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5174;
 end   
18'd167403: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=28;
   mapp<=12;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=4478;
 end   
18'd167404: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=41;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=4841;
 end   
18'd167405: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=30;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=4032;
 end   
18'd167406: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd167407: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd167408: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd167409: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd167410: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd167542: begin  
rid<=1;
end
18'd167543: begin  
end
18'd167544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd167545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd167546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd167547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd167548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd167549: begin  
rid<=0;
end
18'd167601: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=74;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9390;
 end   
18'd167602: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=10;
   mapp<=73;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9075;
 end   
18'd167603: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=19;
   mapp<=78;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=15239;
 end   
18'd167604: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=86;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=15327;
 end   
18'd167605: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=91;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=11421;
 end   
18'd167606: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=4;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=10199;
 end   
18'd167607: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=29;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=13771;
 end   
18'd167608: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=98;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=15966;
 end   
18'd167609: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=48;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd167610: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=37;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd167611: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd167612: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd167613: begin  
  clrr<=0;
  maplen<=3;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9390;
 end   
18'd167742: begin  
rid<=1;
end
18'd167743: begin  
end
18'd167744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd167745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd167746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd167747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd167748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd167749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd167750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd167751: begin  
check<=expctdoutput[7]-outcheck;
end
18'd167752: begin  
rid<=0;
end
18'd167801: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=85;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=24532;
 end   
18'd167802: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=44;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=26796;
 end   
18'd167803: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=83;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd167804: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=6;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd167805: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=11;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd167806: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=7;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd167807: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=6;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd167808: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=82;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd167809: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=92;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd167810: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=8;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd167811: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=94;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd167812: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd167813: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24532;
 end   
18'd167814: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24532;
 end   
18'd167815: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24532;
 end   
18'd167816: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24532;
 end   
18'd167817: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24532;
 end   
18'd167818: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24532;
 end   
18'd167819: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24532;
 end   
18'd167820: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24532;
 end   
18'd167821: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24532;
 end   
18'd167942: begin  
rid<=1;
end
18'd167943: begin  
end
18'd167944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd167945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd167946: begin  
rid<=0;
end
18'd168001: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=43;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=17001;
 end   
18'd168002: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=64;
   mapp<=80;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=21515;
 end   
18'd168003: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=79;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd168004: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=94;
   mapp<=13;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd168005: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=98;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd168006: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd168007: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd168008: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd168009: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd168010: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd168011: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd168142: begin  
rid<=1;
end
18'd168143: begin  
end
18'd168144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd168145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd168146: begin  
rid<=0;
end
18'd168201: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=23;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=253;
 end   
18'd168202: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=34;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=384;
 end   
18'd168203: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=39;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=449;
 end   
18'd168204: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd168342: begin  
rid<=1;
end
18'd168343: begin  
end
18'd168344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd168345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd168346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd168347: begin  
rid<=0;
end
18'd168401: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=81;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5586;
 end   
18'd168402: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=69;
   mapp<=34;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4972;
 end   
18'd168403: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=32;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=3440;
 end   
18'd168404: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=12;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=3141;
 end   
18'd168405: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=31;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=9313;
 end   
18'd168406: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd168407: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd168408: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd168542: begin  
rid<=1;
end
18'd168543: begin  
end
18'd168544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd168545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd168546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd168547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd168548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd168549: begin  
rid<=0;
end
18'd168601: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=82;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=26653;
 end   
18'd168602: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=33;
   mapp<=79;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=32373;
 end   
18'd168603: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=73;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=26294;
 end   
18'd168604: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=95;
   mapp<=69;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=28941;
 end   
18'd168605: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=99;
   mapp<=98;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=24303;
 end   
18'd168606: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=93;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd168607: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd168608: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd168609: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd168610: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd168611: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd168612: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd168613: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26653;
 end   
18'd168614: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26653;
 end   
18'd168615: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26653;
 end   
18'd168616: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26653;
 end   
18'd168742: begin  
rid<=1;
end
18'd168743: begin  
end
18'd168744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd168745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd168746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd168747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd168748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd168749: begin  
rid<=0;
end
18'd168801: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=28;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8567;
 end   
18'd168802: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=86;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6424;
 end   
18'd168803: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=53;
   mapp<=11;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6754;
 end   
18'd168804: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=42;
   mapp<=16;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=11858;
 end   
18'd168805: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=62;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=13697;
 end   
18'd168806: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=42;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=17273;
 end   
18'd168807: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=91;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=16459;
 end   
18'd168808: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd168809: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd168810: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd168811: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd168812: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd168813: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8567;
 end   
18'd168814: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8567;
 end   
18'd168942: begin  
rid<=1;
end
18'd168943: begin  
end
18'd168944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd168945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd168946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd168947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd168948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd168949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd168950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd168951: begin  
rid<=0;
end
18'd169001: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=24;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5004;
 end   
18'd169002: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=81;
   mapp<=52;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5803;
 end   
18'd169003: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=60;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd169004: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd169005: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd169142: begin  
rid<=1;
end
18'd169143: begin  
end
18'd169144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd169145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd169146: begin  
rid<=0;
end
18'd169201: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=76;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3572;
 end   
18'd169202: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=73;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=5558;
 end   
18'd169203: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=59;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=4504;
 end   
18'd169204: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=62;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=4742;
 end   
18'd169205: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=18;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=1408;
 end   
18'd169206: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=54;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=4154;
 end   
18'd169207: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=52;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=4012;
 end   
18'd169208: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=43;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=3338;
 end   
18'd169209: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=4;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=384;
 end   
18'd169210: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd169342: begin  
rid<=1;
end
18'd169343: begin  
end
18'd169344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd169345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd169346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd169347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd169348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd169349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd169350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd169351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd169352: begin  
check<=expctdoutput[8]-outcheck;
end
18'd169353: begin  
rid<=0;
end
18'd169401: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=47;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4371;
 end   
18'd169402: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=9;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=847;
 end   
18'd169403: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd169542: begin  
rid<=1;
end
18'd169543: begin  
end
18'd169544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd169545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd169546: begin  
rid<=0;
end
18'd169601: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=47;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8521;
 end   
18'd169602: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=65;
   mapp<=52;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=14603;
 end   
18'd169603: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=88;
   mapp<=0;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=13453;
 end   
18'd169604: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=4;
   mapp<=1;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=3930;
 end   
18'd169605: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=4;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd169606: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=40;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd169607: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=77;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd169608: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=51;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd169609: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=3;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd169610: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd169611: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd169612: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd169613: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8521;
 end   
18'd169614: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8521;
 end   
18'd169615: begin  
  clrr<=0;
  maplen<=6;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8521;
 end   
18'd169742: begin  
rid<=1;
end
18'd169743: begin  
end
18'd169744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd169745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd169746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd169747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd169748: begin  
rid<=0;
end
18'd169801: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=58;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6701;
 end   
18'd169802: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=15;
   mapp<=85;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7131;
 end   
18'd169803: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=62;
   mapp<=8;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=11426;
 end   
18'd169804: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=72;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=6912;
 end   
18'd169805: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=2;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=6548;
 end   
18'd169806: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=74;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=6898;
 end   
18'd169807: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=6;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=1264;
 end   
18'd169808: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=6;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd169809: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd169810: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd169811: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd169812: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd169942: begin  
rid<=1;
end
18'd169943: begin  
end
18'd169944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd169945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd169946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd169947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd169948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd169949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd169950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd169951: begin  
rid<=0;
end
18'd170001: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=70;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8533;
 end   
18'd170002: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=49;
   mapp<=87;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9579;
 end   
18'd170003: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=71;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=9302;
 end   
18'd170004: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=88;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=7709;
 end   
18'd170005: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=31;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=2700;
 end   
18'd170006: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd170007: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd170008: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd170142: begin  
rid<=1;
end
18'd170143: begin  
end
18'd170144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd170145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd170146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd170147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd170148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd170149: begin  
rid<=0;
end
18'd170201: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=75;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7050;
 end   
18'd170202: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=4;
   mapp<=99;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=14651;
 end   
18'd170203: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=59;
   mapp<=30;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8437;
 end   
18'd170204: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=27;
   mapp<=94;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=13927;
 end   
18'd170205: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=81;
   mapp<=16;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=12256;
 end   
18'd170206: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=20;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd170207: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=38;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd170208: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=83;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd170209: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=10;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd170210: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd170211: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd170212: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd170213: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7050;
 end   
18'd170214: begin  
  clrr<=0;
  maplen<=5;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7050;
 end   
18'd170342: begin  
rid<=1;
end
18'd170343: begin  
end
18'd170344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd170345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd170346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd170347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd170348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd170349: begin  
rid<=0;
end
18'd170401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=15;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4000;
 end   
18'd170402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=59;
   mapp<=40;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5554;
 end   
18'd170403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=40;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd170404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=79;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd170405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd170406: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd170407: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd170542: begin  
rid<=1;
end
18'd170543: begin  
end
18'd170544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd170545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd170546: begin  
rid<=0;
end
18'd170601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=26;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11583;
 end   
18'd170602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=68;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9930;
 end   
18'd170603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=17;
   mapp<=11;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=11650;
 end   
18'd170604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=70;
   mapp<=40;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=8082;
 end   
18'd170605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=15;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd170606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=43;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd170607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd170608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=22;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd170609: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=52;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd170610: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=5;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd170611: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd170612: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd170613: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11583;
 end   
18'd170614: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11583;
 end   
18'd170615: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11583;
 end   
18'd170616: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11583;
 end   
18'd170617: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11583;
 end   
18'd170742: begin  
rid<=1;
end
18'd170743: begin  
end
18'd170744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd170745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd170746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd170747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd170748: begin  
rid<=0;
end
18'd170801: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=16;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10873;
 end   
18'd170802: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=35;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9209;
 end   
18'd170803: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=4;
   mapp<=45;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5280;
 end   
18'd170804: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=18;
   mapp<=40;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=9505;
 end   
18'd170805: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=13;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd170806: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=8;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd170807: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=94;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd170808: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd170809: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd170810: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd170811: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd170812: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd170813: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10873;
 end   
18'd170814: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10873;
 end   
18'd170815: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10873;
 end   
18'd170816: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10873;
 end   
18'd170817: begin  
  clrr<=0;
  maplen<=10;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10873;
 end   
18'd170942: begin  
rid<=1;
end
18'd170943: begin  
end
18'd170944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd170945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd170946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd170947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd170948: begin  
rid<=0;
end
18'd171001: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=81;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6971;
 end   
18'd171002: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=11;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6057;
 end   
18'd171003: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=55;
   mapp<=52;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8115;
 end   
18'd171004: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=48;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=8329;
 end   
18'd171005: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=61;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=6444;
 end   
18'd171006: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=68;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=9551;
 end   
18'd171007: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=13;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=6778;
 end   
18'd171008: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=70;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=9414;
 end   
18'd171009: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd171010: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd171011: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd171012: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd171013: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6971;
 end   
18'd171142: begin  
rid<=1;
end
18'd171143: begin  
end
18'd171144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd171145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd171146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd171147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd171148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd171149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd171150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd171151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd171152: begin  
rid<=0;
end
18'd171201: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=87;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4556;
 end   
18'd171202: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=94;
   mapp<=17;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9103;
 end   
18'd171203: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=81;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=9135;
 end   
18'd171204: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=22;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=10592;
 end   
18'd171205: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=92;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=9360;
 end   
18'd171206: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=14;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=8130;
 end   
18'd171207: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=73;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=8667;
 end   
18'd171208: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=24;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=11276;
 end   
18'd171209: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd171210: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd171211: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd171342: begin  
rid<=1;
end
18'd171343: begin  
end
18'd171344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd171345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd171346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd171347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd171348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd171349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd171350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd171351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd171352: begin  
rid<=0;
end
18'd171401: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=29;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13941;
 end   
18'd171402: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=48;
   mapp<=94;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13143;
 end   
18'd171403: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=53;
   mapp<=29;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12282;
 end   
18'd171404: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=68;
   mapp<=41;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=13094;
 end   
18'd171405: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=58;
   mapp<=81;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=13193;
 end   
18'd171406: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd171407: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd171408: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd171409: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd171410: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd171411: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd171412: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd171413: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13941;
 end   
18'd171414: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13941;
 end   
18'd171542: begin  
rid<=1;
end
18'd171543: begin  
end
18'd171544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd171545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd171546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd171547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd171548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd171549: begin  
rid<=0;
end
18'd171601: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=35;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6556;
 end   
18'd171602: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=78;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd171603: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=13;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd171604: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=44;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd171605: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=59;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd171606: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=16;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd171607: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=2;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd171608: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=13;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd171609: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd171610: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd171611: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd171612: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd171613: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6556;
 end   
18'd171614: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6556;
 end   
18'd171615: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6556;
 end   
18'd171616: begin  
  clrr<=0;
  maplen<=8;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6556;
 end   
18'd171742: begin  
rid<=1;
end
18'd171743: begin  
end
18'd171744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd171745: begin  
rid<=0;
end
18'd171801: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=66;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10607;
 end   
18'd171802: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=18;
   mapp<=27;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11443;
 end   
18'd171803: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=79;
   mapp<=5;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=11859;
 end   
18'd171804: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=43;
   mapp<=24;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=17220;
 end   
18'd171805: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=76;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd171806: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd171807: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd171808: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd171809: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd171810: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd171811: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd171812: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd171813: begin  
  clrr<=0;
  maplen<=8;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10607;
 end   
18'd171942: begin  
rid<=1;
end
18'd171943: begin  
end
18'd171944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd171945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd171946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd171947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd171948: begin  
rid<=0;
end
18'd172001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=34;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16040;
 end   
18'd172002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=22;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd172003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=98;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd172004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=50;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd172005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=46;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd172006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd172007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd172008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd172009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd172010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd172142: begin  
rid<=1;
end
18'd172143: begin  
end
18'd172144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd172145: begin  
rid<=0;
end
18'd172201: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=63;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13892;
 end   
18'd172202: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=64;
   mapp<=46;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11650;
 end   
18'd172203: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=95;
   mapp<=98;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=14508;
 end   
18'd172204: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=26;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=10993;
 end   
18'd172205: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd172206: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd172207: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd172208: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd172209: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd172342: begin  
rid<=1;
end
18'd172343: begin  
end
18'd172344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd172345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd172346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd172347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd172348: begin  
rid<=0;
end
18'd172401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=74;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5566;
 end   
18'd172402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=54;
   mapp<=7;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7051;
 end   
18'd172403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=41;
   mapp<=76;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9937;
 end   
18'd172404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=59;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=6510;
 end   
18'd172405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=27;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=3681;
 end   
18'd172406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=16;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=2506;
 end   
18'd172407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=19;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=5480;
 end   
18'd172408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=6;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=7711;
 end   
18'd172409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=90;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=11827;
 end   
18'd172410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd172411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd172412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd172413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5566;
 end   
18'd172414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5566;
 end   
18'd172542: begin  
rid<=1;
end
18'd172543: begin  
end
18'd172544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd172545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd172546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd172547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd172548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd172549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd172550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd172551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd172552: begin  
check<=expctdoutput[8]-outcheck;
end
18'd172553: begin  
rid<=0;
end
18'd172601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=58;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16750;
 end   
18'd172602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=16;
   mapp<=17;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13358;
 end   
18'd172603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=12;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd172604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=51;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd172605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=71;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd172606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=52;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd172607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd172608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd172609: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd172610: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd172611: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd172612: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd172613: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16750;
 end   
18'd172742: begin  
rid<=1;
end
18'd172743: begin  
end
18'd172744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd172745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd172746: begin  
rid<=0;
end
18'd172801: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=45;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10277;
 end   
18'd172802: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=71;
   mapp<=75;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11628;
 end   
18'd172803: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=62;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd172804: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=45;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd172805: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd172806: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd172807: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd172942: begin  
rid<=1;
end
18'd172943: begin  
end
18'd172944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd172945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd172946: begin  
rid<=0;
end
18'd173001: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=19;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1767;
 end   
18'd173002: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=98;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=1872;
 end   
18'd173003: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=30;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=590;
 end   
18'd173004: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=69;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=1341;
 end   
18'd173005: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=59;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=1161;
 end   
18'd173006: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=73;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=1437;
 end   
18'd173007: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=20;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=440;
 end   
18'd173008: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=85;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=1685;
 end   
18'd173009: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=75;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=1505;
 end   
18'd173010: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=78;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[9]<=1572;
 end   
18'd173011: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd173142: begin  
rid<=1;
end
18'd173143: begin  
end
18'd173144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd173145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd173146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd173147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd173148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd173149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd173150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd173151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd173152: begin  
check<=expctdoutput[8]-outcheck;
end
18'd173153: begin  
check<=expctdoutput[9]-outcheck;
end
18'd173154: begin  
rid<=0;
end
18'd173201: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=79;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=31754;
 end   
18'd173202: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=98;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=30145;
 end   
18'd173203: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=57;
   mapp<=56;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=23824;
 end   
18'd173204: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=69;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd173205: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=45;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd173206: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=48;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd173207: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=65;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd173208: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=67;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd173209: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=21;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd173210: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd173211: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd173212: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd173213: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=31754;
 end   
18'd173214: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=31754;
 end   
18'd173215: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=31754;
 end   
18'd173216: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=31754;
 end   
18'd173342: begin  
rid<=1;
end
18'd173343: begin  
end
18'd173344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd173345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd173346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd173347: begin  
rid<=0;
end
18'd173401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=6;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13542;
 end   
18'd173402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=68;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=14914;
 end   
18'd173403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=92;
   mapp<=32;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=18646;
 end   
18'd173404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=50;
   mapp<=85;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=19412;
 end   
18'd173405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=87;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=19032;
 end   
18'd173406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=93;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=14094;
 end   
18'd173407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=88;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=10738;
 end   
18'd173408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=81;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=12346;
 end   
18'd173409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd173410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=91;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd173411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd173412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd173413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13542;
 end   
18'd173414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13542;
 end   
18'd173415: begin  
  clrr<=0;
  maplen<=11;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13542;
 end   
18'd173542: begin  
rid<=1;
end
18'd173543: begin  
end
18'd173544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd173545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd173546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd173547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd173548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd173549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd173550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd173551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd173552: begin  
rid<=0;
end
18'd173601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=66;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=19474;
 end   
18'd173602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=90;
   mapp<=22;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=19855;
 end   
18'd173603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=39;
   mapp<=34;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=16291;
 end   
18'd173604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=18;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd173605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=65;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd173606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=21;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd173607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=69;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd173608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=89;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd173609: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=58;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd173610: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd173611: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd173612: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd173613: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19474;
 end   
18'd173614: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19474;
 end   
18'd173615: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19474;
 end   
18'd173616: begin  
  clrr<=0;
  maplen<=7;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19474;
 end   
18'd173742: begin  
rid<=1;
end
18'd173743: begin  
end
18'd173744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd173745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd173746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd173747: begin  
rid<=0;
end
18'd173801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=63;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9272;
 end   
18'd173802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=90;
   mapp<=4;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=17477;
 end   
18'd173803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=1;
   mapp<=90;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12770;
 end   
18'd173804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=29;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd173805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=29;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd173806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=47;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd173807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=87;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd173808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=31;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd173809: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd173810: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd173811: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd173812: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd173813: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9272;
 end   
18'd173814: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9272;
 end   
18'd173942: begin  
rid<=1;
end
18'd173943: begin  
end
18'd173944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd173945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd173946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd173947: begin  
rid<=0;
end
18'd174001: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=74;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7500;
 end   
18'd174002: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=40;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9840;
 end   
18'd174003: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=7960;
 end   
18'd174004: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=69;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=6016;
 end   
18'd174005: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=22;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=3228;
 end   
18'd174006: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=39;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=6736;
 end   
18'd174007: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=95;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=9650;
 end   
18'd174008: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd174009: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd174010: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd174142: begin  
rid<=1;
end
18'd174143: begin  
end
18'd174144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd174145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd174146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd174147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd174148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd174149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd174150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd174151: begin  
rid<=0;
end
18'd174201: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=98;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9664;
 end   
18'd174202: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=18;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6750;
 end   
18'd174203: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=6;
   mapp<=5;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=996;
 end   
18'd174204: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=14;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=2632;
 end   
18'd174205: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=39;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=5836;
 end   
18'd174206: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=88;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=10312;
 end   
18'd174207: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd174208: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd174209: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd174210: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd174211: begin  
  clrr<=0;
  maplen<=8;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd174342: begin  
rid<=1;
end
18'd174343: begin  
end
18'd174344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd174345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd174346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd174347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd174348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd174349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd174350: begin  
rid<=0;
end
18'd174401: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=56;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11520;
 end   
18'd174402: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=32;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd174403: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=99;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd174404: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=5;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd174405: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=94;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd174406: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=25;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd174407: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=74;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd174408: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd174409: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd174410: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd174411: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd174412: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd174413: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11520;
 end   
18'd174414: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11520;
 end   
18'd174542: begin  
rid<=1;
end
18'd174543: begin  
end
18'd174544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd174545: begin  
rid<=0;
end
18'd174601: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=47;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=29645;
 end   
18'd174602: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=23;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=29101;
 end   
18'd174603: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=36;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd174604: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=72;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd174605: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=38;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd174606: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=4;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd174607: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=62;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd174608: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=81;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd174609: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=68;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd174610: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=79;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd174611: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd174612: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd174613: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29645;
 end   
18'd174614: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29645;
 end   
18'd174615: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29645;
 end   
18'd174616: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29645;
 end   
18'd174617: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29645;
 end   
18'd174618: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29645;
 end   
18'd174619: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29645;
 end   
18'd174620: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29645;
 end   
18'd174621: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=29645;
 end   
18'd174742: begin  
rid<=1;
end
18'd174743: begin  
end
18'd174744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd174745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd174746: begin  
rid<=0;
end
18'd174801: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=60;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10809;
 end   
18'd174802: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=77;
   mapp<=37;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10035;
 end   
18'd174803: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=27;
   mapp<=30;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12677;
 end   
18'd174804: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=57;
   mapp<=91;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=14932;
 end   
18'd174805: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=7;
   mapp<=49;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=11199;
 end   
18'd174806: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=35;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=12424;
 end   
18'd174807: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=76;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=15394;
 end   
18'd174808: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd174809: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd174810: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd174811: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd174812: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd174813: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10809;
 end   
18'd174814: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10809;
 end   
18'd174815: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10809;
 end   
18'd174816: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10809;
 end   
18'd174942: begin  
rid<=1;
end
18'd174943: begin  
end
18'd174944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd174945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd174946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd174947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd174948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd174949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd174950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd174951: begin  
rid<=0;
end
18'd175001: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=62;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4166;
 end   
18'd175002: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=48;
   mapp<=8;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2946;
 end   
18'd175003: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=1;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=817;
 end   
18'd175004: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=92;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=6346;
 end   
18'd175005: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=88;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=5512;
 end   
18'd175006: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=13;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=987;
 end   
18'd175007: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=18;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=1550;
 end   
18'd175008: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=49;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=3115;
 end   
18'd175009: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=7;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=923;
 end   
18'd175010: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=52;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[9]<=3358;
 end   
18'd175011: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd175012: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd175013: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=4166;
 end   
18'd175142: begin  
rid<=1;
end
18'd175143: begin  
end
18'd175144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd175145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd175146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd175147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd175148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd175149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd175150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd175151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd175152: begin  
check<=expctdoutput[8]-outcheck;
end
18'd175153: begin  
check<=expctdoutput[9]-outcheck;
end
18'd175154: begin  
rid<=0;
end
18'd175201: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=14;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14379;
 end   
18'd175202: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=56;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd175203: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=15;
   mapp<=19;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd175204: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=44;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd175205: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=63;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd175206: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=51;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd175207: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=86;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd175208: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd175209: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd175210: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd175211: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd175212: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd175213: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14379;
 end   
18'd175214: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14379;
 end   
18'd175342: begin  
rid<=1;
end
18'd175343: begin  
end
18'd175344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd175345: begin  
rid<=0;
end
18'd175401: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=81;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=21529;
 end   
18'd175402: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=94;
   mapp<=90;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=14858;
 end   
18'd175403: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=57;
   mapp<=56;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=18831;
 end   
18'd175404: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=72;
   mapp<=59;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=13370;
 end   
18'd175405: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=71;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd175406: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=17;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd175407: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=94;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd175408: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=4;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd175409: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd175410: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd175411: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd175412: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd175413: begin  
  clrr<=0;
  maplen<=5;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21529;
 end   
18'd175542: begin  
rid<=1;
end
18'd175543: begin  
end
18'd175544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd175545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd175546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd175547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd175548: begin  
rid<=0;
end
18'd175601: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=36;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6844;
 end   
18'd175602: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=26;
   mapp<=36;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8770;
 end   
18'd175603: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=52;
   mapp<=70;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6206;
 end   
18'd175604: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=75;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=11023;
 end   
18'd175605: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=3;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=6827;
 end   
18'd175606: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd175607: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=49;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd175608: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd175609: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd175610: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd175742: begin  
rid<=1;
end
18'd175743: begin  
end
18'd175744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd175745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd175746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd175747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd175748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd175749: begin  
rid<=0;
end
18'd175801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=85;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6507;
 end   
18'd175802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=61;
   mapp<=37;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9072;
 end   
18'd175803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=97;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=10217;
 end   
18'd175804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=32;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=5373;
 end   
18'd175805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=43;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=8819;
 end   
18'd175806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd175807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd175808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd175942: begin  
rid<=1;
end
18'd175943: begin  
end
18'd175944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd175945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd175946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd175947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd175948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd175949: begin  
rid<=0;
end
18'd176001: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=4;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=224;
 end   
18'd176002: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=10;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=570;
 end   
18'd176003: begin  
  clrr<=0;
  maplen<=1;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd176142: begin  
rid<=1;
end
18'd176143: begin  
end
18'd176144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd176145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd176146: begin  
rid<=0;
end
18'd176201: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=93;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6672;
 end   
18'd176202: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=75;
   mapp<=22;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7906;
 end   
18'd176203: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=78;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=10799;
 end   
18'd176204: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=47;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=4626;
 end   
18'd176205: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=3;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=7744;
 end   
18'd176206: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=99;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=11282;
 end   
18'd176207: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=27;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=5196;
 end   
18'd176208: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=35;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=9025;
 end   
18'd176209: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd176210: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd176211: begin  
  clrr<=0;
  maplen<=9;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd176342: begin  
rid<=1;
end
18'd176343: begin  
end
18'd176344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd176345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd176346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd176347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd176348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd176349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd176350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd176351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd176352: begin  
rid<=0;
end
18'd176401: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=99;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8710;
 end   
18'd176402: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=14;
   mapp<=14;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1508;
 end   
18'd176403: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=21;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=2736;
 end   
18'd176404: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=65;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd176405: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd176406: begin  
  clrr<=0;
  maplen<=2;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd176542: begin  
rid<=1;
end
18'd176543: begin  
end
18'd176544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd176545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd176546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd176547: begin  
rid<=0;
end
18'd176601: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=25;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4816;
 end   
18'd176602: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=2;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd176603: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=8;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd176604: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd176605: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=33;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd176606: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd176607: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd176608: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd176609: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd176610: begin  
  clrr<=0;
  maplen<=5;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd176742: begin  
rid<=1;
end
18'd176743: begin  
end
18'd176744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd176745: begin  
rid<=0;
end
18'd176801: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=25;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4990;
 end   
18'd176802: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=37;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3347;
 end   
18'd176803: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=26;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=966;
 end   
18'd176804: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=8;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=3190;
 end   
18'd176805: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=80;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=5000;
 end   
18'd176806: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=80;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=5084;
 end   
18'd176807: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=82;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=4219;
 end   
18'd176808: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=57;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=2605;
 end   
18'd176809: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=30;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=4456;
 end   
18'd176810: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd176811: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd176812: begin  
  clrr<=0;
  maplen<=10;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd176942: begin  
rid<=1;
end
18'd176943: begin  
end
18'd176944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd176945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd176946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd176947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd176948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd176949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd176950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd176951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd176952: begin  
check<=expctdoutput[8]-outcheck;
end
18'd176953: begin  
rid<=0;
end
18'd177001: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=69;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5224;
 end   
18'd177002: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=61;
   mapp<=37;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8480;
 end   
18'd177003: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=97;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=8421;
 end   
18'd177004: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=28;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=5439;
 end   
18'd177005: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=57;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=7633;
 end   
18'd177006: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=60;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=5166;
 end   
18'd177007: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd177008: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd177009: begin  
  clrr<=0;
  maplen<=7;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd177142: begin  
rid<=1;
end
18'd177143: begin  
end
18'd177144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd177145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd177146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd177147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd177148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd177149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd177150: begin  
rid<=0;
end
18'd177201: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=4;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=0;
 end   
18'd177202: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=278;
 end   
18'd177203: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=34;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=156;
 end   
18'd177204: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=6;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=54;
 end   
18'd177205: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=92;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=408;
 end   
18'd177206: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=2;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=58;
 end   
18'd177207: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=85;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=400;
 end   
18'd177208: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=16;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=134;
 end   
18'd177209: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=50;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=280;
 end   
18'd177210: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=67;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[9]<=358;
 end   
18'd177211: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=25;
   pp<=100;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[10]<=200;
 end   
18'd177212: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd177342: begin  
rid<=1;
end
18'd177343: begin  
end
18'd177344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd177345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd177346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd177347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd177348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd177349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd177350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd177351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd177352: begin  
check<=expctdoutput[8]-outcheck;
end
18'd177353: begin  
check<=expctdoutput[9]-outcheck;
end
18'd177354: begin  
check<=expctdoutput[10]-outcheck;
end
18'd177355: begin  
rid<=0;
end
18'd177401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=71;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8722;
 end   
18'd177402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=6;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6432;
 end   
18'd177403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=76;
   mapp<=90;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=7235;
 end   
18'd177404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=5;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=5753;
 end   
18'd177405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=59;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=8804;
 end   
18'd177406: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=12;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=14718;
 end   
18'd177407: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=74;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd177408: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=97;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd177409: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd177410: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd177411: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd177542: begin  
rid<=1;
end
18'd177543: begin  
end
18'd177544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd177545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd177546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd177547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd177548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd177549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd177550: begin  
rid<=0;
end
18'd177601: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=80;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14916;
 end   
18'd177602: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=30;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13099;
 end   
18'd177603: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=7;
   mapp<=10;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=16464;
 end   
18'd177604: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=19;
   mapp<=84;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=16054;
 end   
18'd177605: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=13;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd177606: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=74;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd177607: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=55;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd177608: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=32;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd177609: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=92;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd177610: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=56;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd177611: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd177612: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd177613: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14916;
 end   
18'd177614: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14916;
 end   
18'd177615: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14916;
 end   
18'd177616: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14916;
 end   
18'd177617: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14916;
 end   
18'd177742: begin  
rid<=1;
end
18'd177743: begin  
end
18'd177744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd177745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd177746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd177747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd177748: begin  
rid<=0;
end
18'd177801: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=6;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=336;
 end   
18'd177802: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=84;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=514;
 end   
18'd177803: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=2;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=32;
 end   
18'd177804: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=75;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=480;
 end   
18'd177805: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd177942: begin  
rid<=1;
end
18'd177943: begin  
end
18'd177944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd177945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd177946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd177947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd177948: begin  
rid<=0;
end
18'd178001: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=81;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=18974;
 end   
18'd178002: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=58;
   mapp<=54;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=18617;
 end   
18'd178003: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=49;
   mapp<=55;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=18092;
 end   
18'd178004: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=15;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd178005: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=45;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd178006: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=97;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd178007: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=61;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd178008: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=84;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd178009: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd178010: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=25;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd178011: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=62;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd178012: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd178013: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18974;
 end   
18'd178014: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18974;
 end   
18'd178015: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18974;
 end   
18'd178016: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18974;
 end   
18'd178017: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18974;
 end   
18'd178018: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18974;
 end   
18'd178019: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18974;
 end   
18'd178020: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=18974;
 end   
18'd178142: begin  
rid<=1;
end
18'd178143: begin  
end
18'd178144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd178145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd178146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd178147: begin  
rid<=0;
end
18'd178201: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=59;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7224;
 end   
18'd178202: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=4;
   mapp<=50;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5496;
 end   
18'd178203: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=16;
   mapp<=72;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6908;
 end   
18'd178204: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=22;
   mapp<=47;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=4397;
 end   
18'd178205: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=68;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=4650;
 end   
18'd178206: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=62;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=3848;
 end   
18'd178207: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=15;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=2065;
 end   
18'd178208: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd178209: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd178210: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd178211: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd178212: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd178213: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7224;
 end   
18'd178214: begin  
  clrr<=0;
  maplen<=10;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7224;
 end   
18'd178342: begin  
rid<=1;
end
18'd178343: begin  
end
18'd178344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd178345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd178346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd178347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd178348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd178349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd178350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd178351: begin  
rid<=0;
end
18'd178401: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=31;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=961;
 end   
18'd178402: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=3;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=103;
 end   
18'd178403: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=15;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=485;
 end   
18'd178404: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=59;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=1859;
 end   
18'd178405: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=81;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=2551;
 end   
18'd178406: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd178542: begin  
rid<=1;
end
18'd178543: begin  
end
18'd178544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd178545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd178546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd178547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd178548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd178549: begin  
rid<=0;
end
18'd178601: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=72;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=24311;
 end   
18'd178602: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=82;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=24056;
 end   
18'd178603: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=56;
   mapp<=97;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=23593;
 end   
18'd178604: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=82;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd178605: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=93;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd178606: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=47;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd178607: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=55;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd178608: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd178609: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd178610: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd178611: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd178612: begin  
  clrr<=0;
  maplen<=5;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd178742: begin  
rid<=1;
end
18'd178743: begin  
end
18'd178744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd178745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd178746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd178747: begin  
rid<=0;
end
18'd178801: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=7;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=434;
 end   
18'd178802: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=4;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=258;
 end   
18'd178803: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=74;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=4608;
 end   
18'd178804: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd178942: begin  
rid<=1;
end
18'd178943: begin  
end
18'd178944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd178945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd178946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd178947: begin  
rid<=0;
end
18'd179001: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=8;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14068;
 end   
18'd179002: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=63;
   mapp<=9;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=15809;
 end   
18'd179003: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=46;
   mapp<=19;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=18428;
 end   
18'd179004: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=50;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd179005: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=47;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd179006: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=38;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd179007: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=34;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd179008: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd179009: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd179010: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd179011: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd179012: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd179013: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14068;
 end   
18'd179014: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14068;
 end   
18'd179015: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14068;
 end   
18'd179016: begin  
  clrr<=0;
  maplen<=9;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14068;
 end   
18'd179142: begin  
rid<=1;
end
18'd179143: begin  
end
18'd179144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd179145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd179146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd179147: begin  
rid<=0;
end
18'd179201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=59;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6442;
 end   
18'd179202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=80;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=12732;
 end   
18'd179203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=34;
   mapp<=84;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=4614;
 end   
18'd179204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=98;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=10161;
 end   
18'd179205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=27;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd179206: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=56;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd179207: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd179208: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd179209: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd179342: begin  
rid<=1;
end
18'd179343: begin  
end
18'd179344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd179345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd179346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd179347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd179348: begin  
rid<=0;
end
18'd179401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=93;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15101;
 end   
18'd179402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=63;
   mapp<=83;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11671;
 end   
18'd179403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=18;
   mapp<=44;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=11440;
 end   
18'd179404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=61;
   mapp<=65;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=11543;
 end   
18'd179405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=7639;
 end   
18'd179406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd179407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd179408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd179409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd179410: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd179411: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd179412: begin  
  clrr<=0;
  maplen<=8;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd179542: begin  
rid<=1;
end
18'd179543: begin  
end
18'd179544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd179545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd179546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd179547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd179548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd179549: begin  
rid<=0;
end
18'd179601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=67;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5927;
 end   
18'd179602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=93;
   mapp<=8;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5260;
 end   
18'd179603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=4;
   mapp<=48;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=7369;
 end   
18'd179604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=22;
   mapp<=35;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=3392;
 end   
18'd179605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=5;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=4690;
 end   
18'd179606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=39;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=4603;
 end   
18'd179607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd179608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd179609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd179610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd179611: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd179612: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd179613: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5927;
 end   
18'd179742: begin  
rid<=1;
end
18'd179743: begin  
end
18'd179744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd179745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd179746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd179747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd179748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd179749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd179750: begin  
rid<=0;
end
18'd179801: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=79;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=79;
 end   
18'd179802: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=22;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=1748;
 end   
18'd179803: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=9;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=731;
 end   
18'd179804: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=10;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=820;
 end   
18'd179805: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd179942: begin  
rid<=1;
end
18'd179943: begin  
end
18'd179944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd179945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd179946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd179947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd179948: begin  
rid<=0;
end
18'd180001: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=30;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10899;
 end   
18'd180002: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=50;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13262;
 end   
18'd180003: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=49;
   mapp<=83;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=11122;
 end   
18'd180004: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=23;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd180005: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=63;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd180006: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=17;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd180007: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=26;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd180008: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd180009: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd180010: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd180011: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd180012: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd180013: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10899;
 end   
18'd180014: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10899;
 end   
18'd180142: begin  
rid<=1;
end
18'd180143: begin  
end
18'd180144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd180145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd180146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd180147: begin  
rid<=0;
end
18'd180201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=7;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7299;
 end   
18'd180202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=62;
   mapp<=94;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8495;
 end   
18'd180203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=26;
   mapp<=45;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=11833;
 end   
18'd180204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=75;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=12579;
 end   
18'd180205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=81;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=10200;
 end   
18'd180206: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=38;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=12310;
 end   
18'd180207: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=69;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=15635;
 end   
18'd180208: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=92;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd180209: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd180210: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd180211: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd180212: begin  
  clrr<=0;
  maplen<=3;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd180342: begin  
rid<=1;
end
18'd180343: begin  
end
18'd180344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd180345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd180346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd180347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd180348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd180349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd180350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd180351: begin  
rid<=0;
end
18'd180401: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=71;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4488;
 end   
18'd180402: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=9;
   mapp<=49;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4128;
 end   
18'd180403: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=25;
   mapp<=71;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=7286;
 end   
18'd180404: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd180405: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd180406: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd180407: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd180408: begin  
  clrr<=0;
  maplen<=5;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd180542: begin  
rid<=1;
end
18'd180543: begin  
end
18'd180544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd180545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd180546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd180547: begin  
rid<=0;
end
18'd180601: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=1;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10181;
 end   
18'd180602: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=2;
   mapp<=78;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3999;
 end   
18'd180603: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=73;
   mapp<=61;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=10399;
 end   
18'd180604: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=75;
   mapp<=26;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=12278;
 end   
18'd180605: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=3;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd180606: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=24;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd180607: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=29;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd180608: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=49;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd180609: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd180610: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd180611: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd180612: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd180613: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10181;
 end   
18'd180614: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10181;
 end   
18'd180615: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10181;
 end   
18'd180616: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10181;
 end   
18'd180617: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10181;
 end   
18'd180618: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10181;
 end   
18'd180619: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10181;
 end   
18'd180742: begin  
rid<=1;
end
18'd180743: begin  
end
18'd180744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd180745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd180746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd180747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd180748: begin  
rid<=0;
end
18'd180801: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=16;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3711;
 end   
18'd180802: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=47;
   mapp<=49;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3849;
 end   
18'd180803: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=65;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=4632;
 end   
18'd180804: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=76;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=4113;
 end   
18'd180805: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=61;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=5528;
 end   
18'd180806: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=96;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=1727;
 end   
18'd180807: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=3;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=2364;
 end   
18'd180808: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd180809: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd180810: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd180942: begin  
rid<=1;
end
18'd180943: begin  
end
18'd180944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd180945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd180946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd180947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd180948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd180949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd180950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd180951: begin  
rid<=0;
end
18'd181001: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=91;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6993;
 end   
18'd181002: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=59;
   mapp<=74;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3027;
 end   
18'd181003: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=5;
   mapp<=34;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5407;
 end   
18'd181004: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=31;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=9447;
 end   
18'd181005: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=87;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=7493;
 end   
18'd181006: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=63;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=2883;
 end   
18'd181007: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=13;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd181008: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=5;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd181009: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd181010: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd181011: begin  
  clrr<=0;
  maplen<=3;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd181142: begin  
rid<=1;
end
18'd181143: begin  
end
18'd181144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd181145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd181146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd181147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd181148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd181149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd181150: begin  
rid<=0;
end
18'd181201: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=95;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=31632;
 end   
18'd181202: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=23;
   mapp<=51;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=23984;
 end   
18'd181203: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=80;
   mapp<=98;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=24985;
 end   
18'd181204: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=16;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd181205: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=11;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd181206: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=66;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd181207: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=48;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd181208: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=31;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd181209: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd181210: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd181211: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd181212: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd181213: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=31632;
 end   
18'd181214: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=31632;
 end   
18'd181215: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=31632;
 end   
18'd181216: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=31632;
 end   
18'd181217: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=31632;
 end   
18'd181218: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=31632;
 end   
18'd181342: begin  
rid<=1;
end
18'd181343: begin  
end
18'd181344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd181345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd181346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd181347: begin  
rid<=0;
end
18'd181401: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=73;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6321;
 end   
18'd181402: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=53;
   mapp<=38;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3251;
 end   
18'd181403: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=3;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=3883;
 end   
18'd181404: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=97;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=9477;
 end   
18'd181405: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=98;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=8748;
 end   
18'd181406: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=77;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=5581;
 end   
18'd181407: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=26;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd181408: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd181409: begin  
  clrr<=0;
  maplen<=2;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd181542: begin  
rid<=1;
end
18'd181543: begin  
end
18'd181544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd181545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd181546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd181547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd181548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd181549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd181550: begin  
rid<=0;
end
18'd181601: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=69;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=21924;
 end   
18'd181602: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=55;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd181603: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=16;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd181604: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=3;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd181605: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=12;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd181606: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=74;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd181607: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=32;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd181608: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=26;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd181609: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=53;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd181610: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=20;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd181611: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=74;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd181612: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd181613: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21924;
 end   
18'd181614: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21924;
 end   
18'd181615: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21924;
 end   
18'd181616: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21924;
 end   
18'd181617: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21924;
 end   
18'd181618: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21924;
 end   
18'd181619: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21924;
 end   
18'd181620: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21924;
 end   
18'd181621: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21924;
 end   
18'd181622: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=21924;
 end   
18'd181742: begin  
rid<=1;
end
18'd181743: begin  
end
18'd181744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd181745: begin  
rid<=0;
end
18'd181801: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=91;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5070;
 end   
18'd181802: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=91;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2298;
 end   
18'd181803: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=65;
   mapp<=8;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=3127;
 end   
18'd181804: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=24;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=3007;
 end   
18'd181805: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=3;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=6046;
 end   
18'd181806: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=8;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=9540;
 end   
18'd181807: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=77;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=14464;
 end   
18'd181808: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=27;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=10808;
 end   
18'd181809: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd181810: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd181811: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd181812: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd181813: begin  
  clrr<=0;
  maplen<=10;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5070;
 end   
18'd181942: begin  
rid<=1;
end
18'd181943: begin  
end
18'd181944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd181945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd181946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd181947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd181948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd181949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd181950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd181951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd181952: begin  
rid<=0;
end
18'd182001: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=20;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13014;
 end   
18'd182002: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=9;
   mapp<=46;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=12675;
 end   
18'd182003: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=40;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd182004: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=99;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd182005: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=63;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd182006: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=11;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd182007: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=25;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd182008: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=98;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd182009: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=40;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd182010: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=86;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd182011: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd182012: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd182013: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13014;
 end   
18'd182014: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13014;
 end   
18'd182015: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13014;
 end   
18'd182016: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13014;
 end   
18'd182017: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13014;
 end   
18'd182018: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13014;
 end   
18'd182019: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13014;
 end   
18'd182142: begin  
rid<=1;
end
18'd182143: begin  
end
18'd182144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd182145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd182146: begin  
rid<=0;
end
18'd182201: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=52;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5148;
 end   
18'd182202: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=27;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=1414;
 end   
18'd182203: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=73;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=3816;
 end   
18'd182204: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=4;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=238;
 end   
18'd182205: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=76;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=3992;
 end   
18'd182206: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=44;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=2338;
 end   
18'd182207: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=15;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=840;
 end   
18'd182208: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=94;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=4958;
 end   
18'd182209: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=96;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=5072;
 end   
18'd182210: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=13;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[9]<=766;
 end   
18'd182211: begin  
  clrr<=0;
  maplen<=10;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd182342: begin  
rid<=1;
end
18'd182343: begin  
end
18'd182344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd182345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd182346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd182347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd182348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd182349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd182350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd182351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd182352: begin  
check<=expctdoutput[8]-outcheck;
end
18'd182353: begin  
check<=expctdoutput[9]-outcheck;
end
18'd182354: begin  
rid<=0;
end
18'd182401: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=79;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2528;
 end   
18'd182402: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=1;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=89;
 end   
18'd182403: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=31;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=2469;
 end   
18'd182404: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=77;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=6113;
 end   
18'd182405: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=12;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=988;
 end   
18'd182406: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=46;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=3684;
 end   
18'd182407: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=29;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=2351;
 end   
18'd182408: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=67;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=5363;
 end   
18'd182409: begin  
  clrr<=0;
  maplen<=8;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd182542: begin  
rid<=1;
end
18'd182543: begin  
end
18'd182544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd182545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd182546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd182547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd182548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd182549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd182550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd182551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd182552: begin  
rid<=0;
end
18'd182601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=82;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10458;
 end   
18'd182602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=71;
   mapp<=4;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=14337;
 end   
18'd182603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=37;
   mapp<=80;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=15233;
 end   
18'd182604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=70;
   mapp<=4;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=16198;
 end   
18'd182605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=64;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd182606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=65;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd182607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd182608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd182609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd182610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd182611: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd182612: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd182613: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10458;
 end   
18'd182614: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10458;
 end   
18'd182615: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=10458;
 end   
18'd182742: begin  
rid<=1;
end
18'd182743: begin  
end
18'd182744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd182745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd182746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd182747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd182748: begin  
rid<=0;
end
18'd182801: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=25;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=19828;
 end   
18'd182802: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=97;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10922;
 end   
18'd182803: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=10;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=20511;
 end   
18'd182804: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=51;
   mapp<=95;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=10688;
 end   
18'd182805: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=60;
   mapp<=5;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=10716;
 end   
18'd182806: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=62;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd182807: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd182808: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd182809: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd182810: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd182811: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd182812: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd182813: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19828;
 end   
18'd182814: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19828;
 end   
18'd182815: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19828;
 end   
18'd182816: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19828;
 end   
18'd182942: begin  
rid<=1;
end
18'd182943: begin  
end
18'd182944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd182945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd182946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd182947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd182948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd182949: begin  
rid<=0;
end
18'd183001: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=10;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11553;
 end   
18'd183002: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=61;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9981;
 end   
18'd183003: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=78;
   mapp<=81;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5900;
 end   
18'd183004: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=47;
   mapp<=60;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=3675;
 end   
18'd183005: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd183006: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd183007: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd183008: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd183009: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd183010: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd183011: begin  
  clrr<=0;
  maplen<=7;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd183142: begin  
rid<=1;
end
18'd183143: begin  
end
18'd183144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd183145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd183146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd183147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd183148: begin  
rid<=0;
end
18'd183201: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=20;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=25360;
 end   
18'd183202: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=37;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd183203: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=42;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd183204: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=52;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd183205: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=82;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd183206: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=78;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd183207: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=25;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd183208: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=96;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd183209: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=89;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd183210: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=97;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd183211: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=70;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd183212: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd183213: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25360;
 end   
18'd183214: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25360;
 end   
18'd183215: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25360;
 end   
18'd183216: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25360;
 end   
18'd183217: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25360;
 end   
18'd183218: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25360;
 end   
18'd183219: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25360;
 end   
18'd183220: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25360;
 end   
18'd183221: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25360;
 end   
18'd183222: begin  
  clrr<=0;
  maplen<=11;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=25360;
 end   
18'd183342: begin  
rid<=1;
end
18'd183343: begin  
end
18'd183344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd183345: begin  
rid<=0;
end
18'd183401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=86;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15533;
 end   
18'd183402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=69;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=16396;
 end   
18'd183403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=93;
   mapp<=23;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=22749;
 end   
18'd183404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=24;
   mapp<=5;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=23279;
 end   
18'd183405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=60;
   mapp<=72;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=30132;
 end   
18'd183406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=59;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd183407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=95;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd183408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd183409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd183410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd183411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd183412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd183413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15533;
 end   
18'd183414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15533;
 end   
18'd183415: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15533;
 end   
18'd183416: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15533;
 end   
18'd183417: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15533;
 end   
18'd183418: begin  
  clrr<=0;
  maplen<=11;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15533;
 end   
18'd183542: begin  
rid<=1;
end
18'd183543: begin  
end
18'd183544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd183545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd183546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd183547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd183548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd183549: begin  
rid<=0;
end
18'd183601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=3;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=22925;
 end   
18'd183602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=51;
   mapp<=67;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=19675;
 end   
18'd183603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=76;
   mapp<=76;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=17098;
 end   
18'd183604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=42;
   mapp<=2;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=25847;
 end   
18'd183605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=50;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd183606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=98;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd183607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd183608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd183609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd183610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd183611: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd183612: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd183613: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22925;
 end   
18'd183614: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22925;
 end   
18'd183615: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22925;
 end   
18'd183742: begin  
rid<=1;
end
18'd183743: begin  
end
18'd183744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd183745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd183746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd183747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd183748: begin  
rid<=0;
end
18'd183801: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=23;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15534;
 end   
18'd183802: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=78;
   mapp<=56;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=17537;
 end   
18'd183803: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=37;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd183804: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=45;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd183805: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=93;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd183806: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=44;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd183807: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd183808: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd183809: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd183810: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd183811: begin  
  clrr<=0;
  maplen<=5;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd183942: begin  
rid<=1;
end
18'd183943: begin  
end
18'd183944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd183945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd183946: begin  
rid<=0;
end
18'd184001: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=87;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7830;
 end   
18'd184002: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=8;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=730;
 end   
18'd184003: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=85;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=7670;
 end   
18'd184004: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=42;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=3810;
 end   
18'd184005: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=17;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=1570;
 end   
18'd184006: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=19;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=1760;
 end   
18'd184007: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=82;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=7440;
 end   
18'd184008: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=71;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=6460;
 end   
18'd184009: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=30;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=2780;
 end   
18'd184010: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=77;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[9]<=7020;
 end   
18'd184011: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=72;
   mapp<=0;
   pp<=100;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[10]<=6580;
 end   
18'd184012: begin  
  clrr<=0;
  maplen<=1;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd184142: begin  
rid<=1;
end
18'd184143: begin  
end
18'd184144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd184145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd184146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd184147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd184148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd184149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd184150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd184151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd184152: begin  
check<=expctdoutput[8]-outcheck;
end
18'd184153: begin  
check<=expctdoutput[9]-outcheck;
end
18'd184154: begin  
check<=expctdoutput[10]-outcheck;
end
18'd184155: begin  
rid<=0;
end
18'd184201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=46;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5923;
 end   
18'd184202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=35;
   mapp<=45;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6720;
 end   
18'd184203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=29;
   mapp<=50;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=7227;
 end   
18'd184204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=64;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=11262;
 end   
18'd184205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=50;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=11845;
 end   
18'd184206: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=99;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=11517;
 end   
18'd184207: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=84;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=8607;
 end   
18'd184208: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=29;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=7552;
 end   
18'd184209: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=39;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=8497;
 end   
18'd184210: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=78;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd184211: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=49;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd184212: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd184213: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5923;
 end   
18'd184214: begin  
  clrr<=0;
  maplen<=3;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=5923;
 end   
18'd184342: begin  
rid<=1;
end
18'd184343: begin  
end
18'd184344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd184345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd184346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd184347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd184348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd184349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd184350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd184351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd184352: begin  
check<=expctdoutput[8]-outcheck;
end
18'd184353: begin  
rid<=0;
end
18'd184401: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=38;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9363;
 end   
18'd184402: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=65;
   mapp<=35;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=12903;
 end   
18'd184403: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=11;
   mapp<=40;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12723;
 end   
18'd184404: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=73;
   mapp<=64;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=11229;
 end   
18'd184405: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=97;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=14303;
 end   
18'd184406: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=89;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=13619;
 end   
18'd184407: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=7;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd184408: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=91;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd184409: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=79;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd184410: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd184411: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd184412: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd184413: begin  
  clrr<=0;
  maplen<=4;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9363;
 end   
18'd184542: begin  
rid<=1;
end
18'd184543: begin  
end
18'd184544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd184545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd184546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd184547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd184548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd184549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd184550: begin  
rid<=0;
end
18'd184601: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=58;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12921;
 end   
18'd184602: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=17;
   mapp<=49;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=18190;
 end   
18'd184603: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=35;
   mapp<=72;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=14947;
 end   
18'd184604: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=8;
   mapp<=80;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd184605: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=69;
   mapp<=43;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd184606: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=14;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd184607: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=20;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd184608: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=90;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd184609: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=51;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd184610: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd184611: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd184612: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd184613: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12921;
 end   
18'd184614: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12921;
 end   
18'd184615: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12921;
 end   
18'd184616: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12921;
 end   
18'd184617: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12921;
 end   
18'd184618: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12921;
 end   
18'd184619: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12921;
 end   
18'd184620: begin  
  clrr<=0;
  maplen<=11;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12921;
 end   
18'd184742: begin  
rid<=1;
end
18'd184743: begin  
end
18'd184744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd184745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd184746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd184747: begin  
rid<=0;
end
18'd184801: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=15;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5781;
 end   
18'd184802: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=43;
   mapp<=82;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7628;
 end   
18'd184803: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=77;
   mapp<=25;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=3516;
 end   
18'd184804: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=69;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=8158;
 end   
18'd184805: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=2;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=4676;
 end   
18'd184806: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=91;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=2187;
 end   
18'd184807: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=9;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=7879;
 end   
18'd184808: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd184809: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd184810: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd184811: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd184812: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd184942: begin  
rid<=1;
end
18'd184943: begin  
end
18'd184944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd184945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd184946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd184947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd184948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd184949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd184950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd184951: begin  
rid<=0;
end
18'd185001: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=15;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13019;
 end   
18'd185002: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=25;
   mapp<=93;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13882;
 end   
18'd185003: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=28;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd185004: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=75;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd185005: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=55;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd185006: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=41;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd185007: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=53;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd185008: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=10;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd185009: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd185010: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd185011: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd185012: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd185013: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13019;
 end   
18'd185014: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13019;
 end   
18'd185015: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13019;
 end   
18'd185142: begin  
rid<=1;
end
18'd185143: begin  
end
18'd185144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd185145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd185146: begin  
rid<=0;
end
18'd185201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=5;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6297;
 end   
18'd185202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=92;
   mapp<=66;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4612;
 end   
18'd185203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=7;
   mapp<=0;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1853;
 end   
18'd185204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=23;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=6147;
 end   
18'd185205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=77;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=3703;
 end   
18'd185206: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=3;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd185207: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=97;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd185208: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd185209: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd185210: begin  
  clrr<=0;
  maplen<=3;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd185342: begin  
rid<=1;
end
18'd185343: begin  
end
18'd185344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd185345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd185346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd185347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd185348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd185349: begin  
rid<=0;
end
18'd185401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=2;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=114;
 end   
18'd185402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=74;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=158;
 end   
18'd185403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=12;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=44;
 end   
18'd185404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=30;
 end   
18'd185405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=97;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=234;
 end   
18'd185406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=52;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=154;
 end   
18'd185407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=85;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=230;
 end   
18'd185408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=17;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=104;
 end   
18'd185409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=22;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=124;
 end   
18'd185410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=68;
   pp<=90;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[9]<=226;
 end   
18'd185411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=96;
   pp<=100;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[10]<=292;
 end   
18'd185412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd185542: begin  
rid<=1;
end
18'd185543: begin  
end
18'd185544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd185545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd185546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd185547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd185548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd185549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd185550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd185551: begin  
check<=expctdoutput[7]-outcheck;
end
18'd185552: begin  
check<=expctdoutput[8]-outcheck;
end
18'd185553: begin  
check<=expctdoutput[9]-outcheck;
end
18'd185554: begin  
check<=expctdoutput[10]-outcheck;
end
18'd185555: begin  
rid<=0;
end
18'd185601: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=54;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4698;
 end   
18'd185602: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=11;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=967;
 end   
18'd185603: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=70;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6110;
 end   
18'd185604: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd185742: begin  
rid<=1;
end
18'd185743: begin  
end
18'd185744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd185745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd185746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd185747: begin  
rid<=0;
end
18'd185801: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=69;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2652;
 end   
18'd185802: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=17;
   mapp<=87;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6778;
 end   
18'd185803: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=45;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=4723;
 end   
18'd185804: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=94;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=8063;
 end   
18'd185805: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=91;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=7917;
 end   
18'd185806: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=94;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=7522;
 end   
18'd185807: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=58;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=4912;
 end   
18'd185808: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=50;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd185809: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd185810: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd185942: begin  
rid<=1;
end
18'd185943: begin  
end
18'd185944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd185945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd185946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd185947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd185948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd185949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd185950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd185951: begin  
rid<=0;
end
18'd186001: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=52;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=36079;
 end   
18'd186002: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=17;
   mapp<=68;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=33238;
 end   
18'd186003: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=99;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd186004: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=89;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd186005: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=70;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd186006: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=85;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd186007: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=54;
   mapp<=76;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd186008: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=16;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd186009: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=99;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd186010: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=24;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd186011: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=35;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd186012: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd186013: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=36079;
 end   
18'd186014: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=36079;
 end   
18'd186015: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=36079;
 end   
18'd186016: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=36079;
 end   
18'd186017: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=36079;
 end   
18'd186018: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=36079;
 end   
18'd186019: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=36079;
 end   
18'd186020: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=36079;
 end   
18'd186021: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=36079;
 end   
18'd186142: begin  
rid<=1;
end
18'd186143: begin  
end
18'd186144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd186145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd186146: begin  
rid<=0;
end
18'd186201: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=1;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8132;
 end   
18'd186202: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=14;
   mapp<=52;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9766;
 end   
18'd186203: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=85;
   mapp<=56;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=10283;
 end   
18'd186204: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=31;
   mapp<=13;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=5914;
 end   
18'd186205: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=38;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd186206: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=6;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd186207: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=40;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd186208: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=40;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd186209: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd186210: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=17;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd186211: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd186212: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd186213: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8132;
 end   
18'd186214: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8132;
 end   
18'd186215: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8132;
 end   
18'd186216: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8132;
 end   
18'd186217: begin  
  clrr<=0;
  maplen<=7;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8132;
 end   
18'd186342: begin  
rid<=1;
end
18'd186343: begin  
end
18'd186344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd186345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd186346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd186347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd186348: begin  
rid<=0;
end
18'd186401: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=64;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3776;
 end   
18'd186402: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=68;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4022;
 end   
18'd186403: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=12;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=728;
 end   
18'd186404: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=87;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=5163;
 end   
18'd186405: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=46;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=2754;
 end   
18'd186406: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=74;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=4416;
 end   
18'd186407: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=98;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=5842;
 end   
18'd186408: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd186542: begin  
rid<=1;
end
18'd186543: begin  
end
18'd186544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd186545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd186546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd186547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd186548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd186549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd186550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd186551: begin  
rid<=0;
end
18'd186601: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=51;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9827;
 end   
18'd186602: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=17;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=15761;
 end   
18'd186603: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=62;
   mapp<=14;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=14824;
 end   
18'd186604: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=92;
   mapp<=32;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=19303;
 end   
18'd186605: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=52;
   mapp<=65;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=18933;
 end   
18'd186606: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=52;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=11731;
 end   
18'd186607: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=91;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=12376;
 end   
18'd186608: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd186609: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd186610: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd186611: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd186612: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd186613: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9827;
 end   
18'd186614: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9827;
 end   
18'd186615: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9827;
 end   
18'd186616: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=9827;
 end   
18'd186742: begin  
rid<=1;
end
18'd186743: begin  
end
18'd186744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd186745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd186746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd186747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd186748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd186749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd186750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd186751: begin  
rid<=0;
end
18'd186801: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=13;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7022;
 end   
18'd186802: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=18;
   mapp<=8;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6694;
 end   
18'd186803: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=69;
   mapp<=88;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=7130;
 end   
18'd186804: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=57;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=12228;
 end   
18'd186805: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=27;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd186806: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=96;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd186807: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd186808: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd186809: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd186942: begin  
rid<=1;
end
18'd186943: begin  
end
18'd186944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd186945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd186946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd186947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd186948: begin  
rid<=0;
end
18'd187001: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=6;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12706;
 end   
18'd187002: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=30;
   mapp<=44;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=17402;
 end   
18'd187003: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=49;
   mapp<=74;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=19175;
 end   
18'd187004: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=52;
   mapp<=38;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=20566;
 end   
18'd187005: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=57;
   mapp<=98;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=19369;
 end   
18'd187006: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=84;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=17860;
 end   
18'd187007: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=80;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=18112;
 end   
18'd187008: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=72;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd187009: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=52;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd187010: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=43;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd187011: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=69;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd187012: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd187013: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12706;
 end   
18'd187014: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12706;
 end   
18'd187015: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12706;
 end   
18'd187016: begin  
  clrr<=0;
  maplen<=5;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12706;
 end   
18'd187142: begin  
rid<=1;
end
18'd187143: begin  
end
18'd187144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd187145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd187146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd187147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd187148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd187149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd187150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd187151: begin  
rid<=0;
end
18'd187201: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=25;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=19715;
 end   
18'd187202: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=28;
   mapp<=44;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=22353;
 end   
18'd187203: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=41;
   mapp<=8;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd187204: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=77;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd187205: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=25;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd187206: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=82;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd187207: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=11;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd187208: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=78;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd187209: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=61;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd187210: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=96;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd187211: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd187212: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd187213: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19715;
 end   
18'd187214: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19715;
 end   
18'd187215: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19715;
 end   
18'd187216: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19715;
 end   
18'd187217: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19715;
 end   
18'd187218: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19715;
 end   
18'd187219: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19715;
 end   
18'd187220: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19715;
 end   
18'd187221: begin  
  clrr<=0;
  maplen<=11;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19715;
 end   
18'd187342: begin  
rid<=1;
end
18'd187343: begin  
end
18'd187344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd187345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd187346: begin  
rid<=0;
end
18'd187401: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=6;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=162;
 end   
18'd187402: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=34;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=928;
 end   
18'd187403: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=47;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1289;
 end   
18'd187404: begin  
  clrr<=0;
  maplen<=1;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd187542: begin  
rid<=1;
end
18'd187543: begin  
end
18'd187544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd187545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd187546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd187547: begin  
rid<=0;
end
18'd187601: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=83;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=9281;
 end   
18'd187602: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=46;
   mapp<=52;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=7676;
 end   
18'd187603: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=74;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8762;
 end   
18'd187604: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=50;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=7404;
 end   
18'd187605: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=62;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=9242;
 end   
18'd187606: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=78;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=6888;
 end   
18'd187607: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=7;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=3553;
 end   
18'd187608: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=56;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=7162;
 end   
18'd187609: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=47;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=5177;
 end   
18'd187610: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd187611: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd187612: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd187742: begin  
rid<=1;
end
18'd187743: begin  
end
18'd187744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd187745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd187746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd187747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd187748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd187749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd187750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd187751: begin  
check<=expctdoutput[7]-outcheck;
end
18'd187752: begin  
check<=expctdoutput[8]-outcheck;
end
18'd187753: begin  
rid<=0;
end
18'd187801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=93;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=23936;
 end   
18'd187802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=63;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd187803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=2;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd187804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=69;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd187805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=99;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd187806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=80;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd187807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=89;
   mapp<=70;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd187808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd187809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd187810: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd187811: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd187812: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd187813: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23936;
 end   
18'd187814: begin  
  clrr<=0;
  maplen<=7;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=23936;
 end   
18'd187942: begin  
rid<=1;
end
18'd187943: begin  
end
18'd187944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd187945: begin  
rid<=0;
end
18'd188001: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=61;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8074;
 end   
18'd188002: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=18;
   mapp<=66;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8460;
 end   
18'd188003: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=43;
   mapp<=62;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8678;
 end   
18'd188004: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=37;
   mapp<=58;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=9205;
 end   
18'd188005: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=22;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=7162;
 end   
18'd188006: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=78;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=9632;
 end   
18'd188007: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd188008: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd188009: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd188010: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd188011: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd188012: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd188013: begin  
  clrr<=0;
  maplen<=9;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8074;
 end   
18'd188142: begin  
rid<=1;
end
18'd188143: begin  
end
18'd188144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd188145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd188146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd188147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd188148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd188149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd188150: begin  
rid<=0;
end
18'd188201: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=4;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12402;
 end   
18'd188202: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=99;
   mapp<=6;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=17243;
 end   
18'd188203: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=85;
   mapp<=47;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=16026;
 end   
18'd188204: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=39;
   mapp<=29;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd188205: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=92;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd188206: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=6;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd188207: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=27;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd188208: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=16;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd188209: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd188210: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd188211: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd188212: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd188213: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12402;
 end   
18'd188214: begin  
  clrr<=0;
  maplen<=6;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12402;
 end   
18'd188342: begin  
rid<=1;
end
18'd188343: begin  
end
18'd188344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd188345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd188346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd188347: begin  
rid<=0;
end
18'd188401: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=45;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=765;
 end   
18'd188402: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=94;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=4240;
 end   
18'd188403: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=9;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=425;
 end   
18'd188404: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=78;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=3540;
 end   
18'd188405: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=1;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=85;
 end   
18'd188406: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=49;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=2255;
 end   
18'd188407: begin  
  clrr<=0;
  maplen<=6;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd188542: begin  
rid<=1;
end
18'd188543: begin  
end
18'd188544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd188545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd188546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd188547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd188548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd188549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd188550: begin  
rid<=0;
end
18'd188601: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=65;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7523;
 end   
18'd188602: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=87;
   mapp<=1;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5635;
 end   
18'd188603: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=99;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd188604: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=19;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd188605: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd188606: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd188607: begin  
  clrr<=0;
  maplen<=3;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd188742: begin  
rid<=1;
end
18'd188743: begin  
end
18'd188744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd188745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd188746: begin  
rid<=0;
end
18'd188801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=29;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=3270;
 end   
18'd188802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=33;
   mapp<=78;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5014;
 end   
18'd188803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=54;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8570;
 end   
18'd188804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=93;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=9048;
 end   
18'd188805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=87;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=3766;
 end   
18'd188806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=21;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=7964;
 end   
18'd188807: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=95;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=3744;
 end   
18'd188808: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=18;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=6898;
 end   
18'd188809: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=82;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=4310;
 end   
18'd188810: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=29;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd188811: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd188812: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd188942: begin  
rid<=1;
end
18'd188943: begin  
end
18'd188944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd188945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd188946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd188947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd188948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd188949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd188950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd188951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd188952: begin  
check<=expctdoutput[8]-outcheck;
end
18'd188953: begin  
rid<=0;
end
18'd189001: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=39;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1560;
 end   
18'd189002: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=34;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1370;
 end   
18'd189003: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=67;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=2700;
 end   
18'd189004: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=29;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=1190;
 end   
18'd189005: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=79;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=3200;
 end   
18'd189006: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=75;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=3050;
 end   
18'd189007: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=23;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=980;
 end   
18'd189008: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd189142: begin  
rid<=1;
end
18'd189143: begin  
end
18'd189144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd189145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd189146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd189147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd189148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd189149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd189150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd189151: begin  
rid<=0;
end
18'd189201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=38;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11414;
 end   
18'd189202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=81;
   mapp<=88;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=10374;
 end   
18'd189203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=35;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=10020;
 end   
18'd189204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=85;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd189205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=72;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd189206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd189207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd189208: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd189209: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd189210: begin  
  clrr<=0;
  maplen<=4;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd189342: begin  
rid<=1;
end
18'd189343: begin  
end
18'd189344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd189345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd189346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd189347: begin  
rid<=0;
end
18'd189401: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=73;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10615;
 end   
18'd189402: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=70;
   mapp<=70;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6970;
 end   
18'd189403: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=16;
   mapp<=15;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5863;
 end   
18'd189404: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=50;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=9412;
 end   
18'd189405: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=78;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=8204;
 end   
18'd189406: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=17;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=8427;
 end   
18'd189407: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=80;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=12796;
 end   
18'd189408: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd189409: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd189410: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd189411: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd189412: begin  
  clrr<=0;
  maplen<=9;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd189542: begin  
rid<=1;
end
18'd189543: begin  
end
18'd189544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd189545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd189546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd189547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd189548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd189549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd189550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd189551: begin  
rid<=0;
end
18'd189601: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=54;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14365;
 end   
18'd189602: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=12;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd189603: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=49;
   mapp<=61;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd189604: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=75;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd189605: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd189606: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd189607: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd189608: begin  
  clrr<=0;
  maplen<=4;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd189742: begin  
rid<=1;
end
18'd189743: begin  
end
18'd189744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd189745: begin  
rid<=0;
end
18'd189801: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=57;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=26397;
 end   
18'd189802: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=72;
   mapp<=39;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=23066;
 end   
18'd189803: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=74;
   mapp<=94;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=20785;
 end   
18'd189804: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=58;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd189805: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=83;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd189806: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=4;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd189807: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=60;
   mapp<=52;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd189808: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=16;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd189809: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=23;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd189810: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=88;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd189811: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=77;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd189812: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd189813: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26397;
 end   
18'd189814: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26397;
 end   
18'd189815: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26397;
 end   
18'd189816: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26397;
 end   
18'd189817: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26397;
 end   
18'd189818: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26397;
 end   
18'd189819: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26397;
 end   
18'd189820: begin  
  clrr<=0;
  maplen<=9;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=26397;
 end   
18'd189942: begin  
rid<=1;
end
18'd189943: begin  
end
18'd189944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd189945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd189946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd189947: begin  
rid<=0;
end
18'd190001: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=86;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12396;
 end   
18'd190002: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=18;
   mapp<=30;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6397;
 end   
18'd190003: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=81;
   mapp<=54;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=8048;
 end   
18'd190004: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=35;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=9970;
 end   
18'd190005: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd190006: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd190007: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd190008: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd190009: begin  
  clrr<=0;
  maplen<=6;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd190142: begin  
rid<=1;
end
18'd190143: begin  
end
18'd190144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd190145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd190146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd190147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd190148: begin  
rid<=0;
end
18'd190201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=5;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8812;
 end   
18'd190202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=85;
   mapp<=39;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13567;
 end   
18'd190203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=67;
   mapp<=66;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=15277;
 end   
18'd190204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=15;
   mapp<=53;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=11084;
 end   
18'd190205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=98;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=11238;
 end   
18'd190206: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=84;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=10486;
 end   
18'd190207: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=16;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=6565;
 end   
18'd190208: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=26;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=7187;
 end   
18'd190209: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=64;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd190210: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=7;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd190211: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=51;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd190212: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd190213: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8812;
 end   
18'd190214: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8812;
 end   
18'd190215: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8812;
 end   
18'd190342: begin  
rid<=1;
end
18'd190343: begin  
end
18'd190344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd190345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd190346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd190347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd190348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd190349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd190350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd190351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd190352: begin  
rid<=0;
end
18'd190401: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=84;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13135;
 end   
18'd190402: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=65;
   mapp<=51;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=12857;
 end   
18'd190403: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=92;
   mapp<=20;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=14729;
 end   
18'd190404: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=99;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd190405: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=46;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd190406: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd190407: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd190408: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd190542: begin  
rid<=1;
end
18'd190543: begin  
end
18'd190544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd190545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd190546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd190547: begin  
rid<=0;
end
18'd190601: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=3;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=19567;
 end   
18'd190602: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=54;
   mapp<=59;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=22711;
 end   
18'd190603: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=67;
   mapp<=67;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=21855;
 end   
18'd190604: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=95;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd190605: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=58;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd190606: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=57;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd190607: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=57;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd190608: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=69;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd190609: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=22;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd190610: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=4;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd190611: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd190612: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd190613: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19567;
 end   
18'd190614: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19567;
 end   
18'd190615: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19567;
 end   
18'd190616: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19567;
 end   
18'd190617: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19567;
 end   
18'd190618: begin  
  clrr<=0;
  maplen<=8;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=19567;
 end   
18'd190742: begin  
rid<=1;
end
18'd190743: begin  
end
18'd190744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd190745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd190746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd190747: begin  
rid<=0;
end
18'd190801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=68;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12224;
 end   
18'd190802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=3;
   mapp<=17;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4408;
 end   
18'd190803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=47;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd190804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=14;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd190805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=13;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd190806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=5;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd190807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=44;
   mapp<=24;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd190808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=47;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd190809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd190810: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd190811: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd190812: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd190813: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12224;
 end   
18'd190814: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12224;
 end   
18'd190815: begin  
  clrr<=0;
  maplen<=7;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12224;
 end   
18'd190942: begin  
rid<=1;
end
18'd190943: begin  
end
18'd190944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd190945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd190946: begin  
rid<=0;
end
18'd191001: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=56;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6033;
 end   
18'd191002: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=9;
   mapp<=73;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4467;
 end   
18'd191003: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd191004: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd191005: begin  
  clrr<=0;
  maplen<=3;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd191142: begin  
rid<=1;
end
18'd191143: begin  
end
18'd191144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd191145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd191146: begin  
rid<=0;
end
18'd191201: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=12;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=32514;
 end   
18'd191202: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=94;
   mapp<=75;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=40199;
 end   
18'd191203: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=53;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd191204: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=31;
   mapp<=72;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd191205: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=99;
   mapp<=26;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd191206: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=96;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd191207: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=53;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd191208: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=70;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd191209: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=22;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd191210: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=75;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd191211: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd191212: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd191213: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=32514;
 end   
18'd191214: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=32514;
 end   
18'd191215: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=32514;
 end   
18'd191216: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=32514;
 end   
18'd191217: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=32514;
 end   
18'd191218: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=32514;
 end   
18'd191219: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=32514;
 end   
18'd191342: begin  
rid<=1;
end
18'd191343: begin  
end
18'd191344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd191345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd191346: begin  
rid<=0;
end
18'd191401: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=47;
   mapp<=16;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16658;
 end   
18'd191402: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=19;
   mapp<=19;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=19198;
 end   
18'd191403: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=10;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd191404: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=29;
   mapp<=36;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd191405: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=34;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd191406: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=35;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd191407: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=70;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd191408: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=86;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd191409: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=5;
   mapp<=85;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd191410: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=31;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd191411: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=23;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd191412: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd191413: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16658;
 end   
18'd191414: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16658;
 end   
18'd191415: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16658;
 end   
18'd191416: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16658;
 end   
18'd191417: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16658;
 end   
18'd191418: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16658;
 end   
18'd191419: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16658;
 end   
18'd191420: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16658;
 end   
18'd191421: begin  
  clrr<=0;
  maplen<=10;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16658;
 end   
18'd191542: begin  
rid<=1;
end
18'd191543: begin  
end
18'd191544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd191545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd191546: begin  
rid<=0;
end
18'd191601: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=99;
   mapp<=82;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14278;
 end   
18'd191602: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=64;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd191603: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=3;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd191604: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd191605: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd191606: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd191742: begin  
rid<=1;
end
18'd191743: begin  
end
18'd191744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd191745: begin  
rid<=0;
end
18'd191801: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=51;
   mapp<=79;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4029;
 end   
18'd191802: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=13;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1037;
 end   
18'd191803: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=68;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5392;
 end   
18'd191804: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=12;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=978;
 end   
18'd191805: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=8;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=672;
 end   
18'd191806: begin  
  clrr<=0;
  maplen<=1;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd191942: begin  
rid<=1;
end
18'd191943: begin  
end
18'd191944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd191945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd191946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd191947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd191948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd191949: begin  
rid<=0;
end
18'd192001: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=44;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=22277;
 end   
18'd192002: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=46;
   mapp<=94;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=23934;
 end   
18'd192003: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=94;
   mapp<=96;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=20314;
 end   
18'd192004: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=98;
   mapp<=43;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=15517;
 end   
18'd192005: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=25;
   mapp<=64;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=14185;
 end   
18'd192006: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=89;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd192007: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=47;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd192008: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=39;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd192009: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd192010: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd192011: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd192012: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd192013: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22277;
 end   
18'd192014: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22277;
 end   
18'd192015: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22277;
 end   
18'd192016: begin  
  clrr<=0;
  maplen<=10;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22277;
 end   
18'd192142: begin  
rid<=1;
end
18'd192143: begin  
end
18'd192144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd192145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd192146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd192147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd192148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd192149: begin  
rid<=0;
end
18'd192201: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=94;
   mapp<=86;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=32968;
 end   
18'd192202: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=60;
   mapp<=88;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=35690;
 end   
18'd192203: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=98;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd192204: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=62;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd192205: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=98;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd192206: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=32;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd192207: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=47;
   mapp<=42;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd192208: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=77;
   mapp<=88;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd192209: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=33;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd192210: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=52;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd192211: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd192212: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd192213: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=32968;
 end   
18'd192214: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=32968;
 end   
18'd192215: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=32968;
 end   
18'd192216: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=32968;
 end   
18'd192217: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=32968;
 end   
18'd192218: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=32968;
 end   
18'd192219: begin  
  clrr<=0;
  maplen<=9;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=32968;
 end   
18'd192342: begin  
rid<=1;
end
18'd192343: begin  
end
18'd192344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd192345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd192346: begin  
rid<=0;
end
18'd192401: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=97;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4462;
 end   
18'd192402: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=15;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=700;
 end   
18'd192403: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=34;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1584;
 end   
18'd192404: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=54;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=2514;
 end   
18'd192405: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=11;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=546;
 end   
18'd192406: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=37;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=1752;
 end   
18'd192407: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=78;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=3648;
 end   
18'd192408: begin  
  clrr<=0;
  maplen<=1;
  fillen<=7;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd192542: begin  
rid<=1;
end
18'd192543: begin  
end
18'd192544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd192545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd192546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd192547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd192548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd192549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd192550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd192551: begin  
rid<=0;
end
18'd192601: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=13;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8675;
 end   
18'd192602: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=67;
   mapp<=52;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9469;
 end   
18'd192603: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=68;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd192604: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=37;
   mapp<=95;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd192605: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=0;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd192606: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd192607: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd192608: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd192609: begin  
  clrr<=0;
  maplen<=5;
  fillen<=4;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd192742: begin  
rid<=1;
end
18'd192743: begin  
end
18'd192744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd192745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd192746: begin  
rid<=0;
end
18'd192801: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=7;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8045;
 end   
18'd192802: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=29;
   mapp<=48;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9540;
 end   
18'd192803: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=32;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd192804: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=72;
   mapp<=71;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd192805: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=58;
   mapp<=18;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd192806: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd192807: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd192808: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd192809: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd192810: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd192811: begin  
  clrr<=0;
  maplen<=6;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd192942: begin  
rid<=1;
end
18'd192943: begin  
end
18'd192944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd192945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd192946: begin  
rid<=0;
end
18'd193001: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=79;
   mapp<=87;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10063;
 end   
18'd193002: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=55;
   mapp<=58;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4977;
 end   
18'd193003: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=7;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=5248;
 end   
18'd193004: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=85;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=11365;
 end   
18'd193005: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=84;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=8161;
 end   
18'd193006: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=27;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=4603;
 end   
18'd193007: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=44;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=5791;
 end   
18'd193008: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd193009: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd193010: begin  
  clrr<=0;
  maplen<=8;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd193142: begin  
rid<=1;
end
18'd193143: begin  
end
18'd193144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd193145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd193146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd193147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd193148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd193149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd193150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd193151: begin  
rid<=0;
end
18'd193201: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=6;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=8147;
 end   
18'd193202: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=98;
   mapp<=73;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6005;
 end   
18'd193203: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=13;
   mapp<=51;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5437;
 end   
18'd193204: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=43;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=7830;
 end   
18'd193205: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=69;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=6659;
 end   
18'd193206: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=60;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=3302;
 end   
18'd193207: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=25;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=4764;
 end   
18'd193208: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=34;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=10084;
 end   
18'd193209: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=94;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=5451;
 end   
18'd193210: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd193211: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd193212: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd193213: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8147;
 end   
18'd193214: begin  
  clrr<=0;
  maplen<=11;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=8147;
 end   
18'd193342: begin  
rid<=1;
end
18'd193343: begin  
end
18'd193344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd193345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd193346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd193347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd193348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd193349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd193350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd193351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd193352: begin  
check<=expctdoutput[8]-outcheck;
end
18'd193353: begin  
rid<=0;
end
18'd193401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=85;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=24022;
 end   
18'd193402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=62;
   mapp<=54;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=23152;
 end   
18'd193403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=43;
   mapp<=67;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=22268;
 end   
18'd193404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=98;
   mapp<=89;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=24160;
 end   
18'd193405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=3;
   mapp<=65;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=20081;
 end   
18'd193406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=41;
   mapp<=61;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=16605;
 end   
18'd193407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=98;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd193408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=48;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd193409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=4;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd193410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=44;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd193411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=66;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd193412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd193413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24022;
 end   
18'd193414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24022;
 end   
18'd193415: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24022;
 end   
18'd193416: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24022;
 end   
18'd193417: begin  
  clrr<=0;
  maplen<=11;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24022;
 end   
18'd193542: begin  
rid<=1;
end
18'd193543: begin  
end
18'd193544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd193545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd193546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd193547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd193548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd193549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd193550: begin  
rid<=0;
end
18'd193601: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=15;
   mapp<=94;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=24139;
 end   
18'd193602: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=65;
   mapp<=88;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=25552;
 end   
18'd193603: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=81;
   mapp<=21;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=29034;
 end   
18'd193604: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=81;
   mapp<=89;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=30024;
 end   
18'd193605: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=89;
   mapp<=91;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=30137;
 end   
18'd193606: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd193607: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=90;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd193608: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd193609: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=92;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd193610: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd193611: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd193612: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd193613: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24139;
 end   
18'd193614: begin  
  clrr<=0;
  maplen<=9;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=24139;
 end   
18'd193742: begin  
rid<=1;
end
18'd193743: begin  
end
18'd193744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd193745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd193746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd193747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd193748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd193749: begin  
rid<=0;
end
18'd193801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=85;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=10893;
 end   
18'd193802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=84;
   mapp<=87;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=14899;
 end   
18'd193803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=15;
   mapp<=86;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=10222;
 end   
18'd193804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=18;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=9393;
 end   
18'd193805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=92;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=9243;
 end   
18'd193806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd193807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd193808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd193809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd193810: begin  
  clrr<=0;
  maplen<=7;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd193942: begin  
rid<=1;
end
18'd193943: begin  
end
18'd193944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd193945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd193946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd193947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd193948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd193949: begin  
rid<=0;
end
18'd194001: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=47;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4086;
 end   
18'd194002: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=19;
   mapp<=32;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2376;
 end   
18'd194003: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=30;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5408;
 end   
18'd194004: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=99;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=7644;
 end   
18'd194005: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=9;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=1890;
 end   
18'd194006: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=37;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=4356;
 end   
18'd194007: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=49;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=5062;
 end   
18'd194008: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=43;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=5236;
 end   
18'd194009: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=62;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=6940;
 end   
18'd194010: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=71;
   mapp<=0;
   pp<=90;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[9]<=6912;
 end   
18'd194011: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=49;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd194012: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd194013: begin  
  clrr<=0;
  maplen<=2;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=4086;
 end   
18'd194142: begin  
rid<=1;
end
18'd194143: begin  
end
18'd194144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd194145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd194146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd194147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd194148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd194149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd194150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd194151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd194152: begin  
check<=expctdoutput[8]-outcheck;
end
18'd194153: begin  
check<=expctdoutput[9]-outcheck;
end
18'd194154: begin  
rid<=0;
end
18'd194201: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=42;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2058;
 end   
18'd194202: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=4000;
 end   
18'd194203: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=20;
 end   
18'd194204: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=4;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=198;
 end   
18'd194205: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=12;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=544;
 end   
18'd194206: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=42;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=1814;
 end   
18'd194207: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=24;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=1068;
 end   
18'd194208: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=19;
   pp<=70;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[7]<=868;
 end   
18'd194209: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=13;
   pp<=80;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[8]<=626;
 end   
18'd194210: begin  
  clrr<=0;
  maplen<=9;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd194342: begin  
rid<=1;
end
18'd194343: begin  
end
18'd194344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd194345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd194346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd194347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd194348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd194349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd194350: begin  
check<=expctdoutput[6]-outcheck;
end
18'd194351: begin  
check<=expctdoutput[7]-outcheck;
end
18'd194352: begin  
check<=expctdoutput[8]-outcheck;
end
18'd194353: begin  
rid<=0;
end
18'd194401: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=90;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=12400;
 end   
18'd194402: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=97;
   mapp<=13;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11549;
 end   
18'd194403: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=78;
   mapp<=29;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=10605;
 end   
18'd194404: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=1;
   mapp<=13;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=3547;
 end   
18'd194405: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=4;
   mapp<=32;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=6077;
 end   
18'd194406: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=8;
   mapp<=12;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd194407: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=73;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd194408: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=44;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd194409: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=65;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd194410: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=65;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd194411: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd194412: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd194413: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12400;
 end   
18'd194414: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12400;
 end   
18'd194415: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12400;
 end   
18'd194416: begin  
  clrr<=0;
  maplen<=6;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=12400;
 end   
18'd194542: begin  
rid<=1;
end
18'd194543: begin  
end
18'd194544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd194545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd194546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd194547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd194548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd194549: begin  
rid<=0;
end
18'd194601: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=51;
   mapp<=33;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5531;
 end   
18'd194602: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=52;
   mapp<=74;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd194603: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd194604: begin  
  clrr<=0;
  maplen<=2;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd194742: begin  
rid<=1;
end
18'd194743: begin  
end
18'd194744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd194745: begin  
rid<=0;
end
18'd194801: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=96;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=16676;
 end   
18'd194802: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=59;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=14545;
 end   
18'd194803: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=71;
   mapp<=75;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=18969;
 end   
18'd194804: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=2;
   mapp<=74;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=21458;
 end   
18'd194805: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=14;
   mapp<=83;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd194806: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=58;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd194807: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd194808: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=10;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd194809: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd194810: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd194811: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd194812: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd194813: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16676;
 end   
18'd194814: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16676;
 end   
18'd194815: begin  
  clrr<=0;
  maplen<=9;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=16676;
 end   
18'd194942: begin  
rid<=1;
end
18'd194943: begin  
end
18'd194944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd194945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd194946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd194947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd194948: begin  
rid<=0;
end
18'd195001: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=41;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7398;
 end   
18'd195002: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=60;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=11114;
 end   
18'd195003: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=24;
   mapp<=38;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12648;
 end   
18'd195004: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=20;
   mapp<=96;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=10476;
 end   
18'd195005: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=86;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=15062;
 end   
18'd195006: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=81;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=5748;
 end   
18'd195007: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=11;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=10038;
 end   
18'd195008: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=86;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=3222;
 end   
18'd195009: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=12;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd195010: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=34;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd195011: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=5;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd195012: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd195013: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7398;
 end   
18'd195014: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7398;
 end   
18'd195015: begin  
  clrr<=0;
  maplen<=4;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=7398;
 end   
18'd195142: begin  
rid<=1;
end
18'd195143: begin  
end
18'd195144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd195145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd195146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd195147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd195148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd195149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd195150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd195151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd195152: begin  
rid<=0;
end
18'd195201: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=27;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15803;
 end   
18'd195202: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=2;
   mapp<=44;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=12253;
 end   
18'd195203: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=61;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd195204: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=99;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd195205: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=91;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd195206: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=13;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd195207: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=37;
   mapp<=32;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd195208: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=18;
   mapp<=2;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd195209: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=3;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd195210: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd195211: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd195212: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd195213: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15803;
 end   
18'd195214: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15803;
 end   
18'd195215: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15803;
 end   
18'd195216: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15803;
 end   
18'd195217: begin  
  clrr<=0;
  maplen<=8;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15803;
 end   
18'd195342: begin  
rid<=1;
end
18'd195343: begin  
end
18'd195344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd195345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd195346: begin  
rid<=0;
end
18'd195401: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=79;
   mapp<=99;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7821;
 end   
18'd195402: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=42;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=3328;
 end   
18'd195403: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=15;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=1205;
 end   
18'd195404: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=36;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=2874;
 end   
18'd195405: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=1;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=119;
 end   
18'd195406: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=26;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=2104;
 end   
18'd195407: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=54;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=4326;
 end   
18'd195408: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd195542: begin  
rid<=1;
end
18'd195543: begin  
end
18'd195544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd195545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd195546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd195547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd195548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd195549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd195550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd195551: begin  
rid<=0;
end
18'd195601: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=36;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6552;
 end   
18'd195602: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=64;
   mapp<=99;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5245;
 end   
18'd195603: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=49;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=5759;
 end   
18'd195604: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=55;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=8577;
 end   
18'd195605: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=83;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd195606: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd195607: begin  
  clrr<=0;
  maplen<=2;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd195742: begin  
rid<=1;
end
18'd195743: begin  
end
18'd195744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd195745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd195746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd195747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd195748: begin  
rid<=0;
end
18'd195801: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=70;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6140;
 end   
18'd195802: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=10;
   mapp<=9;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=2971;
 end   
18'd195803: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=19;
   mapp<=20;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=3810;
 end   
18'd195804: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=99;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd195805: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=68;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd195806: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd195807: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd195808: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd195942: begin  
rid<=1;
end
18'd195943: begin  
end
18'd195944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd195945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd195946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd195947: begin  
rid<=0;
end
18'd196001: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=41;
   mapp<=30;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=15883;
 end   
18'd196002: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=81;
   mapp<=18;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=21708;
 end   
18'd196003: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=78;
   mapp<=17;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=16390;
 end   
18'd196004: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=82;
   mapp<=2;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=14687;
 end   
18'd196005: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=7;
   mapp<=77;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd196006: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=97;
   mapp<=34;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd196007: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=90;
   mapp<=68;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd196008: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=76;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd196009: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=33;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd196010: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=21;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd196011: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=80;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd196012: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd196013: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15883;
 end   
18'd196014: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15883;
 end   
18'd196015: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15883;
 end   
18'd196016: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15883;
 end   
18'd196017: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15883;
 end   
18'd196018: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15883;
 end   
18'd196019: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=15883;
 end   
18'd196142: begin  
rid<=1;
end
18'd196143: begin  
end
18'd196144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd196145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd196146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd196147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd196148: begin  
rid<=0;
end
18'd196201: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=87;
   mapp<=41;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11757;
 end   
18'd196202: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=37;
   mapp<=34;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8358;
 end   
18'd196203: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=57;
   mapp<=8;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=14683;
 end   
18'd196204: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=70;
   mapp<=26;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=11133;
 end   
18'd196205: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=20;
   mapp<=39;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=12805;
 end   
18'd196206: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=51;
   mapp<=76;
   pp<=50;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=10211;
 end   
18'd196207: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=24;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd196208: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=99;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd196209: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=35;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd196210: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=80;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd196211: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=32;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd196212: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd196213: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11757;
 end   
18'd196214: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11757;
 end   
18'd196215: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11757;
 end   
18'd196216: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11757;
 end   
18'd196217: begin  
  clrr<=0;
  maplen<=6;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11757;
 end   
18'd196342: begin  
rid<=1;
end
18'd196343: begin  
end
18'd196344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd196345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd196346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd196347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd196348: begin  
check<=expctdoutput[4]-outcheck;
end
18'd196349: begin  
check<=expctdoutput[5]-outcheck;
end
18'd196350: begin  
rid<=0;
end
18'd196401: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=76;
   mapp<=60;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4560;
 end   
18'd196402: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=77;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=5862;
 end   
18'd196403: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=86;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=6556;
 end   
18'd196404: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=17;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=1322;
 end   
18'd196405: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=1;
   pp<=40;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[4]<=116;
 end   
18'd196406: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=46;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=3546;
 end   
18'd196407: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=68;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=5228;
 end   
18'd196408: begin  
  clrr<=0;
  maplen<=7;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd196542: begin  
rid<=1;
end
18'd196543: begin  
end
18'd196544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd196545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd196546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd196547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd196548: begin  
check<=expctdoutput[4]-outcheck;
end
18'd196549: begin  
check<=expctdoutput[5]-outcheck;
end
18'd196550: begin  
check<=expctdoutput[6]-outcheck;
end
18'd196551: begin  
rid<=0;
end
18'd196601: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=88;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=7524;
 end   
18'd196602: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=68;
   mapp<=34;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=9751;
 end   
18'd196603: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=61;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd196604: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=17;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd196605: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd196606: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd196607: begin  
  clrr<=0;
  maplen<=4;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd196742: begin  
rid<=1;
end
18'd196743: begin  
end
18'd196744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd196745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd196746: begin  
rid<=0;
end
18'd196801: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=17;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1529;
 end   
18'd196802: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=32;
   mapp<=9;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1955;
 end   
18'd196803: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=56;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=1164;
 end   
18'd196804: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=6;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd196805: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd196806: begin  
  clrr<=0;
  maplen<=4;
  fillen<=2;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd196942: begin  
rid<=1;
end
18'd196943: begin  
end
18'd196944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd196945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd196946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd196947: begin  
rid<=0;
end
18'd197001: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=11;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2747;
 end   
18'd197002: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=30;
   mapp<=78;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8140;
 end   
18'd197003: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=90;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=9980;
 end   
18'd197004: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=85;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=10819;
 end   
18'd197005: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=98;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=8970;
 end   
18'd197006: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=68;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=5218;
 end   
18'd197007: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=34;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=1396;
 end   
18'd197008: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=1;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=5801;
 end   
18'd197009: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=73;
   mapp<=0;
   pp<=80;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[8]<=5355;
 end   
18'd197010: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=33;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd197011: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd197012: begin  
  clrr<=0;
  maplen<=2;
  fillen<=10;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd197142: begin  
rid<=1;
end
18'd197143: begin  
end
18'd197144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd197145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd197146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd197147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd197148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd197149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd197150: begin  
check<=expctdoutput[6]-outcheck;
end
18'd197151: begin  
check<=expctdoutput[7]-outcheck;
end
18'd197152: begin  
check<=expctdoutput[8]-outcheck;
end
18'd197153: begin  
rid<=0;
end
18'd197201: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=40;
   mapp<=53;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2120;
 end   
18'd197202: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=5;
   pp<=10;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[1]<=210;
 end   
18'd197203: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=20;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[2]<=20;
 end   
18'd197204: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=4;
   pp<=30;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[3]<=190;
 end   
18'd197205: begin  
  clrr<=0;
  maplen<=4;
  fillen<=1;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd197342: begin  
rid<=1;
end
18'd197343: begin  
end
18'd197344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd197345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd197346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd197347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd197348: begin  
rid<=0;
end
18'd197401: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=16;
   mapp<=45;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=13143;
 end   
18'd197402: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=53;
   mapp<=95;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=21451;
 end   
18'd197403: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=93;
   mapp<=22;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=12859;
 end   
18'd197404: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=48;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=19474;
 end   
18'd197405: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=95;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd197406: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=50;
   mapp<=96;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd197407: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=32;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd197408: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=75;
   mapp<=3;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd197409: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=67;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd197410: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=97;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd197411: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=38;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd197412: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd197413: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13143;
 end   
18'd197414: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13143;
 end   
18'd197415: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13143;
 end   
18'd197416: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13143;
 end   
18'd197417: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13143;
 end   
18'd197418: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13143;
 end   
18'd197419: begin  
  clrr<=0;
  maplen<=11;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=13143;
 end   
18'd197542: begin  
rid<=1;
end
18'd197543: begin  
end
18'd197544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd197545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd197546: begin  
check<=expctdoutput[2]-outcheck;
end
18'd197547: begin  
check<=expctdoutput[3]-outcheck;
end
18'd197548: begin  
rid<=0;
end
18'd197601: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=14;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5771;
 end   
18'd197602: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=17;
   mapp<=20;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[1]<=10;
 end   
18'd197603: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=73;
   mapp<=65;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd197604: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd197605: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd197606: begin  
  clrr<=0;
  maplen<=3;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd197742: begin  
rid<=1;
end
18'd197743: begin  
end
18'd197744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd197745: begin  
rid<=0;
end
18'd197801: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=36;
   mapp<=27;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=4104;
 end   
18'd197802: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=58;
   mapp<=54;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6868;
 end   
18'd197803: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=98;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6608;
 end   
18'd197804: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=73;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=4215;
 end   
18'd197805: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=41;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=2389;
 end   
18'd197806: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=23;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=2129;
 end   
18'd197807: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=27;
   mapp<=0;
   pp<=60;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[6]<=5919;
 end   
18'd197808: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=95;
   mapp<=0;
   pp<=70;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[7]<=3121;
 end   
18'd197809: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=9;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd197810: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd197811: begin  
  clrr<=0;
  maplen<=2;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd197942: begin  
rid<=1;
end
18'd197943: begin  
end
18'd197944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd197945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd197946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd197947: begin  
check<=expctdoutput[3]-outcheck;
end
18'd197948: begin  
check<=expctdoutput[4]-outcheck;
end
18'd197949: begin  
check<=expctdoutput[5]-outcheck;
end
18'd197950: begin  
check<=expctdoutput[6]-outcheck;
end
18'd197951: begin  
check<=expctdoutput[7]-outcheck;
end
18'd197952: begin  
rid<=0;
end
18'd198001: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=69;
   mapp<=23;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1587;
 end   
18'd198002: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=64;
   mapp<=0;
   pp<=10;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=1482;
 end   
18'd198003: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=55;
   mapp<=0;
   pp<=20;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=1285;
 end   
18'd198004: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=34;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=812;
 end   
18'd198005: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=95;
   mapp<=0;
   pp<=40;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=2225;
 end   
18'd198006: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=53;
   mapp<=0;
   pp<=50;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[5]<=1269;
 end   
18'd198007: begin  
  clrr<=0;
  maplen<=1;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd198142: begin  
rid<=1;
end
18'd198143: begin  
end
18'd198144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd198145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd198146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd198147: begin  
check<=expctdoutput[3]-outcheck;
end
18'd198148: begin  
check<=expctdoutput[4]-outcheck;
end
18'd198149: begin  
check<=expctdoutput[5]-outcheck;
end
18'd198150: begin  
rid<=0;
end
18'd198201: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=10;
   mapp<=11;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1685;
 end   
18'd198202: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=18;
   mapp<=79;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4309;
 end   
18'd198203: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=51;
   mapp<=3;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=2705;
 end   
18'd198204: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=24;
   mapp<=0;
   pp<=30;
   gm<=0;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=6415;
 end   
18'd198205: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=76;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd198206: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=39;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd198207: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd198208: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd198209: begin  
  clrr<=0;
  maplen<=3;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd198342: begin  
rid<=1;
end
18'd198343: begin  
end
18'd198344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd198345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd198346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd198347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd198348: begin  
rid<=0;
end
18'd198401: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=52;
   mapp<=62;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=5384;
 end   
18'd198402: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=30;
   mapp<=72;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=3382;
 end   
18'd198403: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=21;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd198404: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd198405: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd198542: begin  
rid<=1;
end
18'd198543: begin  
end
18'd198544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd198545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd198546: begin  
rid<=0;
end
18'd198601: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=61;
   mapp<=51;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=14338;
 end   
18'd198602: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=54;
   mapp<=71;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=8146;
 end   
18'd198603: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=2;
   mapp<=11;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=13412;
 end   
18'd198604: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=87;
   mapp<=83;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=9101;
 end   
18'd198605: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=30;
   mapp<=5;
   pp<=40;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[4]<=11582;
 end   
18'd198606: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=87;
   pp<=50;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[5]<=13804;
 end   
18'd198607: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=22;
   pp<=60;
   gm<=1;
   gf<=0;
   gp<=1;
 expctdoutput[6]<=12757;
 end   
18'd198608: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=55;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd198609: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=57;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd198610: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=73;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd198611: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=64;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd198612: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd198613: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14338;
 end   
18'd198614: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14338;
 end   
18'd198615: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14338;
 end   
18'd198616: begin  
  clrr<=0;
  maplen<=11;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=14338;
 end   
18'd198742: begin  
rid<=1;
end
18'd198743: begin  
end
18'd198744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd198745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd198746: begin  
check<=expctdoutput[2]-outcheck;
end
18'd198747: begin  
check<=expctdoutput[3]-outcheck;
end
18'd198748: begin  
check<=expctdoutput[4]-outcheck;
end
18'd198749: begin  
check<=expctdoutput[5]-outcheck;
end
18'd198750: begin  
check<=expctdoutput[6]-outcheck;
end
18'd198751: begin  
rid<=0;
end
18'd198801: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=62;
   mapp<=28;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=6376;
 end   
18'd198802: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=25;
   mapp<=51;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=5134;
 end   
18'd198803: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=7;
   mapp<=14;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd198804: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=43;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd198805: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=79;
   mapp<=0;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd198806: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=6;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd198807: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd198808: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd198809: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd198810: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd198811: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd198812: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd198813: begin  
  clrr<=0;
  maplen<=7;
  fillen<=6;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=6376;
 end   
18'd198942: begin  
rid<=1;
end
18'd198943: begin  
end
18'd198944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd198945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd198946: begin  
rid<=0;
end
18'd199001: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=9;
   mapp<=54;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=2401;
 end   
18'd199002: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=19;
   mapp<=65;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=4246;
 end   
18'd199003: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=34;
   mapp<=20;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=6126;
 end   
18'd199004: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=50;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd199005: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=51;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd199006: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd199007: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd199008: begin  
  clrr<=0;
  maplen<=3;
  fillen<=5;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd199142: begin  
rid<=1;
end
18'd199143: begin  
end
18'd199144: begin  
check<=expctdoutput[0]-outcheck;
end
18'd199145: begin  
check<=expctdoutput[1]-outcheck;
end
18'd199146: begin  
check<=expctdoutput[2]-outcheck;
end
18'd199147: begin  
rid<=0;
end
18'd199201: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=7;
   mapp<=1;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=17313;
 end   
18'd199202: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=3;
   mapp<=38;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=17104;
 end   
18'd199203: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=22;
   mapp<=46;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=20036;
 end   
18'd199204: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=59;
   mapp<=77;
   pp<=30;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[3]<=18713;
 end   
18'd199205: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=15;
   mapp<=58;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd199206: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=59;
   mapp<=81;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd199207: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=55;
   mapp<=49;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd199208: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=89;
   mapp<=37;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd199209: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=4;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd199210: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=52;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd199211: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=83;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd199212: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd199213: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17313;
 end   
18'd199214: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17313;
 end   
18'd199215: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17313;
 end   
18'd199216: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17313;
 end   
18'd199217: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17313;
 end   
18'd199218: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17313;
 end   
18'd199219: begin  
  clrr<=0;
  maplen<=8;
  fillen<=11;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=17313;
 end   
18'd199342: begin  
rid<=1;
end
18'd199343: begin  
end
18'd199344: begin  
check<=expctdoutput[0]-outcheck;
end
18'd199345: begin  
check<=expctdoutput[1]-outcheck;
end
18'd199346: begin  
check<=expctdoutput[2]-outcheck;
end
18'd199347: begin  
check<=expctdoutput[3]-outcheck;
end
18'd199348: begin  
rid<=0;
end
18'd199401: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=4;
   mapp<=93;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=1792;
 end   
18'd199402: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=20;
   mapp<=71;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=6414;
 end   
18'd199403: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=64;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd199404: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd199405: begin  
  clrr<=0;
  maplen<=2;
  fillen<=3;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd199542: begin  
rid<=1;
end
18'd199543: begin  
end
18'd199544: begin  
check<=expctdoutput[0]-outcheck;
end
18'd199545: begin  
check<=expctdoutput[1]-outcheck;
end
18'd199546: begin  
rid<=0;
end
18'd199601: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=95;
   mapp<=25;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=11320;
 end   
18'd199602: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=3;
   mapp<=0;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=13907;
 end   
18'd199603: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=9;
   mapp<=21;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[2]<=20;
 end   
18'd199604: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=6;
   mapp<=78;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd199605: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=92;
   mapp<=7;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd199606: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=83;
   mapp<=31;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd199607: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=31;
   mapp<=35;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd199608: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=22;
   mapp<=59;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd199609: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=48;
   mapp<=56;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd199610: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=89;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd199611: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd199612: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd199613: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11320;
 end   
18'd199614: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11320;
 end   
18'd199615: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11320;
 end   
18'd199616: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11320;
 end   
18'd199617: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11320;
 end   
18'd199618: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11320;
 end   
18'd199619: begin  
  clrr<=0;
  maplen<=10;
  fillen<=9;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=11320;
 end   
18'd199742: begin  
rid<=1;
end
18'd199743: begin  
end
18'd199744: begin  
check<=expctdoutput[0]-outcheck;
end
18'd199745: begin  
check<=expctdoutput[1]-outcheck;
end
18'd199746: begin  
rid<=0;
end
18'd199801: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=56;
   mapp<=15;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[0]<=22434;
 end   
18'd199802: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=36;
   mapp<=28;
   pp<=10;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[1]<=24200;
 end   
18'd199803: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=97;
   mapp<=68;
   pp<=20;
   gm<=1;
   gf<=1;
   gp<=1;
 expctdoutput[2]<=23039;
 end   
18'd199804: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=77;
   mapp<=84;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[3]<=30;
 end   
18'd199805: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=63;
   mapp<=46;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[4]<=40;
 end   
18'd199806: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=38;
   mapp<=63;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[5]<=50;
 end   
18'd199807: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=37;
   mapp<=40;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[6]<=60;
 end   
18'd199808: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=10;
   mapp<=75;
   pp<=0;
   gm<=1;
   gf<=1;
   gp<=0;
 expctdoutput[7]<=70;
 end   
18'd199809: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=22;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[8]<=80;
 end   
18'd199810: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=69;
   pp<=0;
   gm<=1;
   gf<=0;
   gp<=0;
 expctdoutput[9]<=90;
 end   
18'd199811: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[10]<=100;
 end   
18'd199812: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[11]<=110;
 end   
18'd199813: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22434;
 end   
18'd199814: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22434;
 end   
18'd199815: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22434;
 end   
18'd199816: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22434;
 end   
18'd199817: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22434;
 end   
18'd199818: begin  
  clrr<=0;
  maplen<=10;
  fillen<=8;
   filterp<=0;
   mapp<=0;
   pp<=0;
   gm<=0;
   gf<=0;
   gp<=0;
 expctdoutput[0]<=22434;
 end   
18'd199942: begin  
rid<=1;
end
18'd199943: begin  
end
18'd199944: begin  
check<=expctdoutput[0]-outcheck;
end
18'd199945: begin  
check<=expctdoutput[1]-outcheck;
end
18'd199946: begin  
check<=expctdoutput[2]-outcheck;
end
18'd199947: begin  
rid<=0;
end







 endcase

end


endmodule